s, ma'am. What can I get you today?""

""I'd like 12 scotches, neat.""

Thinking that's a bit of an odd order, he pours her a stiff one and sets it on the bar. 

""Slam!"", she downs that drink like a free beer at a Geological Society of America convention. 

""Keep'em coming..."" she purrs.

One after another. 10, 9, 8 and all that. She drains those 11 scotches without so much as a hiccup. She pays up, thanks the barkeep, slumps like a poleaxed mule and passes out colder'n a mackerel. 

The barkeep looks over the bar at her, slumped between the peanut hulls and cigarette butts on the floor. Some of the regulars saunter over and inspect the scene as well. 

""Well"", says Shady (a regular regular), ""What'd we do with her now?""

""Y'know..."", offers Earl (another regular), ""She's so out of it, we could all have a wee bit of the ol' in/out/in/out, and she'd never be the wiser...just sayin'""

A chorus of ""Hell yeah's"" and ""Firsties!"" rebound around the bar.

After the deeds were done, she was cleaned up, her purse inspected, her address ascertained,  a cab called and she was sent on her way home.  

The very next day, she infiltrates the bar again and...

 Confidently saunters up to the bar and hails the barman.

""Yes, ma'am. What can I get you today?""

""I'd like 12 scotches, neat.""

""Coming up.""

A dozen drinks later, the exact same scenario plays out.  The Lagavulin-slam, wipeout, rumpy-pumpy, deshevilization,  cab called, etc.

The very next day, she infiltrates the bar again and...

""Good day, Ma'am."" exclaims the barkeep. ""Your usual?""

""No, not today. Today I'd like 12 vodkas. Those damn scotches make my pussy hurt...""
",This rather attractive woman walks into a bar...,2
post,4q3wps,2qh72,jokes,false,1467041366,https://old.reddit.com/r/Jokes/comments/4q3wps/gay_jokes_arnt_funny/,self.jokes,,Come on guys.,Gay jokes arn't funny,9
post,4q3w37,2qh72,jokes,false,1467041169,https://old.reddit.com/r/Jokes/comments/4q3w37/a_classic_that_my_dad_has_always_told_me_i_am/,self.jokes,,"Roses are red,


Violets are blue,


You have an arranged marriage waiting for you",A classic that my dad has always told me (I am Indian immigrant),0
post,4q3vrz,2qh72,jokes,false,1467041066,https://old.reddit.com/r/Jokes/comments/4q3vrz/how_much_space_had_the_eu_freed/,self.jokes,,[deleted],How much space had the EU freed?,0
post,4q3v3b,2qh72,jokes,false,1467040851,https://old.reddit.com/r/Jokes/comments/4q3v3b/bhola_was_busy_in_removing_a_wheel_from_auto3/,self.jokes,,"ramu:why are you removing a wheel from auto?
bhola:can't you read ""parking for two wheelers only""",Bhola was busy in removing a wheel from auto(3 wheeler)...,1
post,4q3uvk,2qh72,jokes,false,1467040776,https://old.reddit.com/r/Jokes/comments/4q3uvk/make_sure_you_tip_your_waitress/,self.jokes,,It's very funny when they fall over.,Make sure you tip your waitress...,38
post,4q3u1u,2qh72,jokes,false,1467040512,https://old.reddit.com/r/Jokes/comments/4q3u1u/where_was_tommen_found_when_he_jumped_off_the_roof/,self.jokes,,King's landing.,Where was Tommen found when he jumped off the roof?,1
post,4q3txm,2qh72,jokes,false,1467040476,https://old.reddit.com/r/Jokes/comments/4q3txm/vegans/,self.jokes,,Please don't downvote,Vegans,0
post,4q3twv,2qh72,jokes,false,1467040469,https://old.reddit.com/r/Jokes/comments/4q3twv/roses_are_red_violets_are_blue/,self.jokes,,"This poem doesn't rhyme.

Refrigerator ","Roses are red, violets are blue...",0
post,4q3tws,2qh72,jokes,false,1467040467,https://old.reddit.com/r/Jokes/comments/4q3tws/what_is_the_fastest_thing_you_know/,self.jokes,,"""What is the fastest thing you know?""  the interviewer asked to 4 candidates.

Dave, the American, replied,""A THOUGHT”. It just pops into your head. There's no warning that it's on the way; it's just there. A thought is the fastest thing I know of.""

""That's very good!"" replied the interviewer. 
""And now you sir?"" he asked Vladimir , the Russian.

""Hmm... let me see. A blink! It comes and goes and you don't know that it ever happened. A BLINK is the fastest thing I know.

""Excellent!"" said the interviewer. ""The blink of an eye, that's a very popular cliché for speed”. 

He then turned to George, the Australian who was contemplating his reply.

""Well, out at my dad's ranch, you step out of the house and on the wall there's a light switch. When you flip that switch, way out across the pasture the light in the barn comes on. Yep, Turning on a LIGHT is the fastest thing I can think of.""

The interviewer was very impressed with the third answer and thought he had found his man. ""It's hard to beat the speed of light"" he said.

Turning to Patel, the Guy from India , the fourth and final man, the interviewer posed the same question. 

Patel replied, (in his Gujju accent!) ""Apter herring da 3 prebius ansers sir, et's obius to me dat the fastest thing is DIARRHEA.""

""WHAT!?"" said the interviewer, stunned by the response. The others were already giggling in their seats..

""Oh, I can expleyn sir,"" said Patel. “You see, sir, da ader day my tummy was pheeling bad and so I run so fast to the baatrum, but before I could THINK, BLINK, or TURN ON THE LIGHT, I alredi done it !

""Patel is now the new ""Office Manager"" at Wal-Mart in Washington.
","""What is the fastest thing you know?""",95
post,4q3tir,2qh72,jokes,false,1467040361,https://old.reddit.com/r/Jokes/comments/4q3tir/3_friends_are_boasting_about_their_grandfathers/,self.jokes,,"James: Do you know my grandpa's unusual talent? He can drink one liter of water in one breath. Yep, that's how talented he is.


Jeff: You call that a talent? You're grandpa has nothing on mine. Can your grandpa sleep while standing? When my grandpa feels sleepy, he just closes his eyes while standing and instantly falls asleep on the spot; without leaning on any support.


Steven: Your grandpas are such untalented piece of shits. My grandpa brushes his teeth while smoking a cigarette.


Jeff: Is your grandpa retarded? It would be impossible to not get the cigarette wet!


Steven: Oh he does it easily. He removes his dentures first.",3 friends are boasting about their grandfathers' most unusual talents..,0
post,4q3swc,2qh72,jokes,false,1467040161,https://old.reddit.com/r/Jokes/comments/4q3swc/little_audrey/,self.jokes,,"Little Audrey was sitting on the porch with her younger brother when she said, “Look, there’s a quarter in the street!” Her brother jumped up and ran into the street to get the money and was promptly squashed by a truck.

Little Audrey laughed and laughed, because she knew it was only a nickel.",Little Audrey...,6
post,4q3so3,2qh72,jokes,false,1467040086,https://old.reddit.com/r/Jokes/comments/4q3so3/if_the_majority_of_people_in_the_us_celebrate/,self.jokes,,Then the amount of people that celebrate Hanukkah are in the menorahty,If the majority of people in the US celebrate Christmas,3
post,4q3sfv,2qh72,jokes,false,1467040008,https://old.reddit.com/r/Jokes/comments/4q3sfv/comedy_news_6272016/,self.jokes,,"Independence Day weekend is coming up. When we celebrate the courage of our ancestors by grilling fattening food, arguing with relatives and watching drunk uncle Remus blow off a few more fingers! God bless America!

The BET Black Entertainment Awards were held over the weekend. Hey, wasn't it just 5 months ago that the Academy Awards were slammed for not having enough African Americans?

On this  day in 1963 JFK visited Ireland. prompting his famous comment, ""Wow, Don't they ever sober up?""

Donald Trump has come out against gay marriage. He says marriage is a holy &amp; sacred institution between a rich man and his trophy wife.

The stock market is going crazy since the Brexit. It's like an orgy; Pants are down skirts are up &amp; everybody's getting screwed!

Some people still don't believe in climate change despite the fact the term was coined by George Bush. So tell me is Bush a liar, or is it real?

Finding Dory is number one at the box office, It's kind of an animated 'Home Alone' underwater.

A friend invited me to a weekend at a nudist colony. Nudity (if you're not a supermodel or athlete) is something that works better in concept form!

Today's Inspirational Thought; I'm always shocked at how consistently great life can be...if you let it.

The Girl Scouts are allegedly 347 mill in debt. Don't worry, they plan to fix the problem by raising cookie prices to $175. a box!

Scientist claim men are predisposed to looking at other women. And women are predisposed to elbowing men in the ribs as hard as possible!

 I believe this is Gay Pride Week in New York. You can tell by the outrageous clothes, wild makeup &amp; outlandish behavior. No wait...it's New York, that;s normal.

A Racine, Wisconsin man died after taking too big a bite of a piece of meat. It's known as 'Mama Cass Syndrome'. 

",Comedy News 6/27/2016,0
post,4q3ra9,2qh72,jokes,false,1467039651,https://old.reddit.com/r/Jokes/comments/4q3ra9/you_wont_believe_what_they_called_their_online/,self.jokes,,Click Bait,You won't believe what they called their online store for fishing tackle!,1
post,4q3r9d,2qh72,jokes,false,1467039642,https://old.reddit.com/r/Jokes/comments/4q3r9d/a_koala_walks_into_a_bar/,self.jokes,,"So he sits down and after a while of chatting with the barkeep he starts to notice a girl eyeing him from across the bar. So he goes and talks to her and after some flirting they decide to go upstairs

So they go upstairs and get into the 69 position and when its all said and done the koala goes to leave, but the girl says ""Hey, where's my money?"" Appalled he says ""What do you mean?"" She replies by telling him to look up the definition of prostitute in the dictionary. He does so and it reads 'One who does sexual acts for money.' He then tells her to look up the definition of koala in the dictionary. She does this and it reads ""small, tree dwelling marsupial that eats bush and leaves.""",A Koala walks into a bar...,90
post,4q3qwn,2qh72,jokes,false,1467039529,https://old.reddit.com/r/Jokes/comments/4q3qwn/rjokes_flair_system/,self.jokes,,[removed],/r/jokes flair system,1
post,4q3qqr,2qh72,jokes,false,1467039480,https://old.reddit.com/r/Jokes/comments/4q3qqr/its_been_reported_that_donald_trump_has_recently/,self.jokes,,And had him deported. ,It's been reported that Donald Trump has recently found Jesus ...,760
post,4q3q8t,2qh72,jokes,false,1467039328,https://old.reddit.com/r/Jokes/comments/4q3q8t/weather_for_all/,self.jokes,,[removed],Weather for All,1
post,4q3q88,2qh72,jokes,false,1467039321,https://old.reddit.com/r/Jokes/comments/4q3q88/guess_well_be_seeing_more_of_ronaldo_on_the_cover/,self.jokes,,or is the Barstillona ?,Guess we'll be seeing more of Ronaldo on the cover of EA Fifa now..,1
post,4q3pui,2qh72,jokes,false,1467039210,https://old.reddit.com/r/Jokes/comments/4q3pui/how_does_luke_skywalker_masturbate/,self.jokes,,Han Solo ,How does Luke Skywalker masturbate?,0
post,4q3pib,2qh72,jokes,false,1467039095,https://old.reddit.com/r/Jokes/comments/4q3pib/dvds_are_dying_because_of_torrents/,self.jokes,,[deleted],DVDs are dying because of torrents,0
post,4q3p8p,2qh72,jokes,false,1467039006,https://old.reddit.com/r/Jokes/comments/4q3p8p/you_cant_trust_a_mule_with_an_important_task/,self.jokes,,They'll just half-ass it.,You can't trust a mule with an important task.,29
post,4q3ozw,2qh72,jokes,false,1467038917,https://old.reddit.com/r/Jokes/comments/4q3ozw/how_does_pinocchios_father_know_when_his_son/,self.jokes,,He just nose it.,How does Pinocchio's father know when his son tells a lie?,10
post,4q3oko,2qh72,jokes,false,1467038778,https://old.reddit.com/r/Jokes/comments/4q3oko/an_american_an_englishman_and_a_scotsman_walk/,self.jokes,,"They all order a pint of best bitter, when a fly lands in each ones glass. 

The American picks the fly out, and consumes his beer.

The Englishman asks the barman politely for another beer. 

The Scotsman deftly picks the fly out of his beer, and starts slamming it on the rim of the glass howling ""Give it back, ya wee bastard!""","An American, an Englishman and a Scotsman walk into a bar...",4
post,4q3nce,2qh72,jokes,false,1467038376,https://old.reddit.com/r/Jokes/comments/4q3nce/swimming_pool_wishes/,self.jokes,,"    At a swimming pool: Three guys climb a high-dive tower and meet a good fairy who offers to fulfill a wish for each of them. One jumps and says, ""Beer!"" - and the pool is full of beer. The other one jumps, says, ""Money!"" and the pool is full of money. The last one starts to jump but slips and, falling, yells, ""SHIIIIIIT!!!""
",swimming pool wishes,18
post,4q3mx7,2qh72,jokes,false,1467038225,https://old.reddit.com/r/Jokes/comments/4q3mx7/kids_today/,self.jokes,,"I was out at the pub quiz with my nieces and nephews the other night, and the final round was all about Matt Damon films. We got absolutely trounced.

Kids today don't know their Bourne.",Kids today...,0
post,4q3mi5,2qh72,jokes,false,1467038094,https://old.reddit.com/r/Jokes/comments/4q3mi5/a_couple_is_going_through_a_divorce/,self.jokes,,"The mom makes a big fuss, saying she absolutely HAS to keep the son. The dad asks ""Why?""

""Because I gave birth to him!""

The man thinks for a while and finally says ""If I put money into a soda vending machine, is the soda mine or the machine's?""",a couple is going through a divorce,12
post,4q3mi2,2qh72,jokes,false,1467038093,https://old.reddit.com/r/Jokes/comments/4q3mi2/who_speaks_latin/,self.jokes,,[deleted],Who speaks Latin?,0
post,4q3m1b,2qh72,jokes,false,1467037936,https://old.reddit.com/r/Jokes/comments/4q3m1b/why_do_australians_take_forever_to_play_chess/,self.jokes,,"Because they never make it past the first check, mate.",Why do Australians take forever to play chess?,4
post,4q3llw,2qh72,jokes,false,1467037794,https://old.reddit.com/r/Jokes/comments/4q3llw/one_night_a_scottish_couple_took_a_walk_through_a/,self.jokes,,"The woman says to the man, ''You want to hold my hand, don't you?''

The man says,''Yes, how did you know?'' 

She says, ''By the gleam in your eye.'' 

So they held hands. 

A little down the road the woman says to the man, ''You want to kiss me don't you?'' 

The man says,''Yes, how did you know?'' 

She says, ''By the gleam in your eye.'' 

So they kissed and kept walking. 

A little later the woman askes the man, ''You want to screw me don't you?''

 The man says, ''How did you know? By the gleam in my eye?'' 

The woman says, ''No, by the tilt in your kilt.''",One night a Scottish couple took a walk through a beautiful lit up town...,8
post,4q3lk4,2qh72,jokes,false,1467037780,https://old.reddit.com/r/Jokes/comments/4q3lk4/my_dad_has_a_weird_obsession/,self.jokes,,[deleted],My dad has a weird obsession...,0
post,4q3jpk,2qh72,jokes,false,1467037132,https://old.reddit.com/r/Jokes/comments/4q3jpk/you_gotta_love_north_korea/,self.jokes,,[deleted],You gotta love north korea...,919
post,4q3j28,2qh72,jokes,false,1467036907,https://old.reddit.com/r/Jokes/comments/4q3j28/what_is_a_small_update_to_a_guitar_chord_app/,self.jokes,,Am update,What is a small update to a Guitar Chord app called?,0
post,4q3id6,2qh72,jokes,false,1467036645,https://old.reddit.com/r/Jokes/comments/4q3id6/whats_the_best_thing_about_naming_your_dog_rihanna/,self.jokes,,"You know when you beat it, she will keep coming back to you!",What's the best thing about naming your dog Rihanna?,0
post,4q3hod,2qh72,jokes,false,1467036390,https://old.reddit.com/r/Jokes/comments/4q3hod/i_needed_to_upgrade_my_car_sound_system/,self.jokes,,"So I put a gimp suit on my dog and put her in the trunk, now I have a new subwoofer.",I needed to upgrade my car sound system,1
post,4q3heo,2qh72,jokes,false,1467036289,https://old.reddit.com/r/Jokes/comments/4q3heo/i_dont_have_any_idea_how_to_fix_this_hole_in_my/,self.jokes,,Darn it.,I don't have any idea how to fix this hole in my jumper...,0
post,4q3gzd,2qh72,jokes,false,1467036131,https://old.reddit.com/r/Jokes/comments/4q3gzd/to_be_stung_by_a_mosquito_is_not_very_pleasant/,self.jokes,,"But the thought that an insect with just 10 brain cells could mess up your entire night is something quite different.

",To be stung by a mosquito is not very pleasant...,0
post,4q3grf,2qh72,jokes,false,1467036053,https://old.reddit.com/r/Jokes/comments/4q3grf/what_happened_to_the_man_with_a_legal_fetish_when/,self.jokes,,He got off on a technicality,What happened to the man with a legal fetish when he went to court for his parking ticket?,30
post,4q3fqm,2qh72,jokes,false,1467035659,https://old.reddit.com/r/Jokes/comments/4q3fqm/the_news_of_kings_landing_destruction_mustve/,self.jokes,,[removed],The news of Kings Landing destruction must've spread through Westeros like...,0
post,4q3fe9,2qh72,jokes,false,1467035551,https://old.reddit.com/r/Jokes/comments/4q3fe9/have_you_heard_about_the_new_superpopular_broom/,self.jokes,,It's sweeping the nation,Have you heard about the new super-popular broom that came out?,12
post,4q3ent,2qh72,jokes,false,1467035292,https://old.reddit.com/r/Jokes/comments/4q3ent/nsfw_my_new_girlfriend_just_introduced_me_to_her/,self.jokes,,"I didn't want to tell anyone, but I just had to get this shit off my chest.",[NSFW] My new girlfriend just introduced me to her fetish....,212
post,4q3ei6,2qh72,jokes,false,1467035222,https://old.reddit.com/r/Jokes/comments/4q3ei6/what_was_that_justin_timberlake_song_about_the/,self.jokes,,[deleted],What was that Justin Timberlake song about the Chornaya?,2
post,4q3dhu,2qh72,jokes,false,1467034849,https://old.reddit.com/r/Jokes/comments/4q3dhu/why_didnt_the_alcoholic_become_a_lawyer/,self.jokes,,because he couldn't pass the bar,why didn't the alcoholic become a lawyer?,18
post,4q3dhf,2qh72,jokes,false,1467034845,https://old.reddit.com/r/Jokes/comments/4q3dhf/bartender_theres_a_fly_in_my_beer/,self.jokes,,"A millionaire, a hard hat, and an old drunk are at a bar. When they get their beers, they notice a fly in each mug.
The millionaire politely asks the bartender for another beer, then proceeds to sip it.
The hard hat spills out just enough to get rid of the fly and quaffs the rest.
It's now the old drunk's turn. He sticks his hand into the beer, grabs the fly by the wings, and shouts, ""Spit it out! Spit it out!""","Bartender, There's a Fly In My Beer!",7
post,4q3cut,2qh72,jokes,false,1467034605,https://old.reddit.com/r/Jokes/comments/4q3cut/what_does_samuel_l_jackson_say/,self.jokes,,"When you’re about to throw your cigarette in the street?

“Hold on to your butts.”


When you’re bleeding from multiple stab wounds?

“Hold on to your cuts.”


When someone from Holland is forgetting their language?

“Hold on to your dutch.” 


When someone is being eaten by a velociraptor?

“Hold on to your guts.”


When a hurricane is heading towards a South Pacific Island?

“Hold on to your huts.”


When you’re dangling from a cliff?

“Hold on to your juts.”


When you’re adopting dogs from the pound?

“Hold on to your mutts.“


When he’s playing paintball?

“Hold onto your nuts.”


When he’s playing mini-golf?

“Hold on to your putts.” 


When you’re having a bubble bath?

“Hold on to your suds.” 


When he picks his nose?

“Mmm hmm, this is a tasty booger!” 

(edit: thanks pickles)
",What does Samuel L. Jackson say...,0
post,4q3bwh,2qh72,jokes,false,1467034223,https://old.reddit.com/r/Jokes/comments/4q3bwh/three_men_are_standing_in_front_of_the_heavens/,self.jokes,,[deleted],Three men are standing in front of the heavens door,1
post,4q3buo,2qh72,jokes,false,1467034209,https://old.reddit.com/r/Jokes/comments/4q3buo/what_noise_do_the_the_irish_make_when_theyre/,self.jokes,,[deleted],What noise do the the Irish make when they're kicked out of Europe?,1
post,4q3btu,2qh72,jokes,false,1467034197,https://old.reddit.com/r/Jokes/comments/4q3btu/what_do_you_call_a_damaged_instrument_in_the_16th/,self.jokes,,B-roke ,What do you call a damaged instrument in the 16th century?,1
post,4q3ahn,2qh72,jokes,false,1467033706,https://old.reddit.com/r/Jokes/comments/4q3ahn/i_called_my_husband_to_get_something_for_the_kids/,self.jokes,,[deleted],I called my husband to get something for the kids.,0
post,4q397k,2qh72,jokes,false,1467033208,https://old.reddit.com/r/Jokes/comments/4q397k/a_terrorist_is_at_your_door/,self.jokes,,[deleted],A terrorist is at your door.,0
post,4q38y3,2qh72,jokes,false,1467033121,https://old.reddit.com/r/Jokes/comments/4q38y3/do_strangers_shit_in_the_woods/,self.jokes,,"Yes. I happened, incidentally, and quite unfortunately, to turn a corner in a local forest to see a guy shitting in the woods. And I did not turn the soft bend to see his face as he was squeezing, no, I turned and saw his ass.

This was public lands no more than 100 yards from a cafe and beaches where families swim.

HILARIOUS!",Do strangers shit in the woods?,0
post,4q386t,2qh72,jokes,false,1467032829,https://old.reddit.com/r/Jokes/comments/4q386t/a_couple_is_going_through_a_divorce_and_custody/,self.jokes,,"The father presents evidence that the wife hits the poor boy whenever he misbehaves the slightest. The mother reveals evidence that the father would get belligerently drunk and use his belt on the boy.

The Judge suggests letting the boy live with his grandfather, but it turns out that almost everyone in this twisted family has a history of domestic violence. Not wanting to subject the poor boy to a life of physical punishment, the court decided to take a recess to brainstorm what to do with the son. The court eventually comes to a historic and unprecedented conclusion:

The boy would be in custody of the England national football team because they're incapable of beating anyone.   ",A couple is going through a divorce and custody of the son comes into question.,2215
post,4q37xy,2qh72,jokes,false,1467032720,https://old.reddit.com/r/Jokes/comments/4q37xy/little_april_was_not_the_best_student_in_sunday/,self.jokes,,[removed],Little April was not the best student in Sunday school.,1
post,4q37f2,2qh72,jokes,false,1467032502,https://old.reddit.com/r/Jokes/comments/4q37f2/fifa_games/,self.jokes,,[deleted],Fifa Games.,0
post,4q35s6,2qh72,jokes,false,1467031843,https://old.reddit.com/r/Jokes/comments/4q35s6/why_arent_digital_images_of_bob_marley_scalable/,self.jokes,,Because they're all rasta graphics.,Why aren't digital images of Bob Marley scalable?,15
post,4q355h,2qh72,jokes,false,1467031583,https://old.reddit.com/r/Jokes/comments/4q355h/an_englishman_a_scotsman_and_an_irishman_walk/,self.jokes,,"An Englishman, a Scotsman and an Irishman walk into a bar...

The Englishman wanted to go so they all had to leave.","An Englishman, a Scotsman and an Irishman walk into a bar...",17590
post,4q33bg,2qh72,jokes,false,1467030857,https://old.reddit.com/r/Jokes/comments/4q33bg/doctor_patient/,self.jokes,,[deleted],Doctor &amp; Patient,0
post,4q33a4,2qh72,jokes,false,1467030843,https://old.reddit.com/r/Jokes/comments/4q33a4/attention_attention/,self.jokes,,"
Please... "" Lifebuoy "" Do not get bathed ,
.
.
They hear "" Kidao "" ko Maarta Hai ..
.
.
And "" you "" do not want to lose .",** Attention ** ** Attention **,0
post,4q32es,2qh72,jokes,false,1467030488,https://old.reddit.com/r/Jokes/comments/4q32es/i_played_a_blank_cd_full_blast_on_repeat_all/,self.jokes,,The mime next door went nuts!,I played a blank CD full blast on repeat all night last night.,34
post,4q320p,2qh72,jokes,false,1467030323,https://old.reddit.com/r/Jokes/comments/4q320p/if_trump_becomes_president_it_wont_be_called_the/,self.jokes,,He'll rename it the Exclusively White House,"If Trump becomes president, it won't be called the White House anymore",0
post,4q31dl,2qh72,jokes,false,1467030032,https://old.reddit.com/r/Jokes/comments/4q31dl/after_news_of_brexit_australia_is_set_to_leave/,self.jokes,,They would like to be known as just Stralia now.,"After news of Brexit, Australia is set to leave the AU",0
post,4q2znk,2qh72,jokes,false,1467029230,https://old.reddit.com/r/Jokes/comments/4q2znk/nobody_uses_dvds_most_of_em_use_torrents/,self.jokes,,Hence DVD Rip,Nobody uses DVDs. Most of em' use Torrents.,3
post,4q2yqo,2qh72,jokes,false,1467028792,https://old.reddit.com/r/Jokes/comments/4q2yqo/why_did_the_eu_start_downloading_random_stuff_to/,self.jokes,,It had freed up one GB of space.,Why did the EU start downloading random stuff to it's computer?,13
post,4q2y7j,2qh72,jokes,false,1467028544,https://old.reddit.com/r/Jokes/comments/4q2y7j/a_monk_to_another_o_master_is_it_proper_for_a/,self.jokes,,"""Sure, as long as there are no attachments"", replied the other.","A monk to another, ""O! master, is it proper for a monk to use email?""",3
post,4q2y09,2qh72,jokes,false,1467028434,https://old.reddit.com/r/Jokes/comments/4q2y09/a_young_man_is_in_a_terrible_accident/,self.jokes,,"and as a result he loses one of his eyes. 
He goes to see the optician and the Dr says ""I'm sorry sir, but we're all out of new glass eyes, so we can only offer one of the old wooden eyes"".
The young man accepts and leaves the clinic.
That weekend he heads to a local dance, everyone is dancing around and having fun except for one girl all alone, the man's friend spots her and says ""go and ask her for a dance"".
The young man gets up the courage to head over and taps her on the shoulder:
""Excuse me miss, would you like to dance?""
The girl turns around and peculiarly has her mouth vertical instead of horizontal.
She is overjoyed with being asked to dance and exclaims back ""Oh wow, wouldn't I!""
To which the young man yells back, ""Oi, don't call me wooden eye, cunt mouth!""
",A young man is in a terrible accident,7
post,4q2xu5,2qh72,jokes,false,1467028333,https://old.reddit.com/r/Jokes/comments/4q2xu5/why_was_cinderella_kicked_out_of_the_football_team/,self.jokes,,She ran away from the ball.,Why was Cinderella kicked out of the football team?,89
post,4q2xop,2qh72,jokes,false,1467028256,https://old.reddit.com/r/Jokes/comments/4q2xop/jumpoline/,self.jokes,,"They used to call it a Jumpoline, until your mum went on it.",Jumpoline,0
post,4q2xlk,2qh72,jokes,false,1467028215,https://old.reddit.com/r/Jokes/comments/4q2xlk/how_do_you_find_will_smith_in_the_snow/,self.jokes,,You look for fresh prints.,How do you find Will Smith in the snow?,0
post,4q2xce,2qh72,jokes,false,1467028074,https://old.reddit.com/r/Jokes/comments/4q2xce/well_done_to_wales_for_putting_northern_ireland/,self.jokes,,[removed],Well done to Wales for putting Northern Ireland out of Europe twice in one week...,1
post,4q2wrw,2qh72,jokes,false,1467027768,https://old.reddit.com/r/Jokes/comments/4q2wrw/classic_joke_for_our_muslim_friends_today/,self.jokes,,"There were two white christian men, John and Mike, whose plane crashed into a desert. Luckily they survived unharmed. As they traveled through the hot desert looking for food and water, they gave up and sat down, thinking of what to do.

As the dust in the air settled, they suddenly could view a mosque ahead. They became very hopeful. But then John said ''Muslims are there. They might help us if we say we are Muslim.'' Then Mike said ''No way, I won't say I'm Muslim, I'm gonna be honest''.

So John and Mike went to the Mosque ahead and were greeted by an Arab Muslim, who asked what their names were.

John thought of a Muslim name and said, 'My name is Muhammad'. And Mike said 'My name is Mike'.

The Arab man said 'Hello Mike.' And told these other men to take Mike and give him food and drink.

Then he turned to John and said, 'Salaam Muhammad. Ramadan Mubarak! (Hello Muhammad, Happy Ramadan)
",Classic joke for our Muslim friends today,1074
post,4q2wnr,2qh72,jokes,false,1467027716,https://old.reddit.com/r/Jokes/comments/4q2wnr/a_philosopher_a_mathematician_and_an_idiot_were/,self.jokes,,[deleted],"A philosopher, a mathematician and an idiot were riding in a car when it crashed into a tree",0
post,4q2wj7,2qh72,jokes,false,1467027645,https://old.reddit.com/r/Jokes/comments/4q2wj7/so_they_are_making_a_new_ghostbusters_with_a/,self.jokes,,"Apparently it's not going to be called ""Ballbusters""",So they are making a new ghostbusters with a female cast,0
post,4q2w8b,2qh72,jokes,false,1467027500,https://old.reddit.com/r/Jokes/comments/4q2w8b/a_local_prison_introduced_an_english_literature/,self.jokes,,".. during the inmates' free time. The thought behind it was that if the prisoners had lessons on great writers such as Joyce, Hemingway, or Poe it would help them express themselves as well as helping with their rehabilitation back into society. Unfortunately, the program failed. It seems that when choosing where to spend their time, the prisoners preferred the cons to prose.",A local prison introduced an English Literature course...,6
post,4q2vwk,2qh72,jokes,false,1467027327,https://old.reddit.com/r/Jokes/comments/4q2vwk/why_was_iagos_plan_so_well_calculated/,self.jokes,,[deleted],Why was Iago's plan so well calculated?,0
post,4q2vmp,2qh72,jokes,false,1467027178,https://old.reddit.com/r/Jokes/comments/4q2vmp/if_you_find_faith_in_religion_just_remember_it/,self.jokes,,[removed],If you find faith in religion just remember it should be a long term commitment rather than a fad.,0
post,4q2v96,2qh72,jokes,false,1467026973,https://old.reddit.com/r/Jokes/comments/4q2v96/whats_the_difference_between_english_breakfast/,self.jokes,,One is still in the EU.,Whats the difference between English Breakfast and Irish Breakfast tea?,0
post,4q2v23,2qh72,jokes,false,1467026863,https://old.reddit.com/r/Jokes/comments/4q2v23/the_eu_just_formed_a_dance_group/,self.jokes,,"It's called ""free movement""",The EU just formed a dance group!,0
post,4q2u82,2qh72,jokes,false,1467026422,https://old.reddit.com/r/Jokes/comments/4q2u82/why_was_iagos_plans_so_well_calculated/,self.jokes,,[deleted],Why was Iago's plans so well calculated?,1
post,4q2teq,2qh72,jokes,false,1467025958,https://old.reddit.com/r/Jokes/comments/4q2teq/all_that_voted_for_brexit_should_be_jailed_for/,self.jokes,,Because they want to fuck an entire generation of kids.,All that voted for Brexit should be jailed for pedophilia...,0
post,4q2tdu,2qh72,jokes,false,1467025946,https://old.reddit.com/r/Jokes/comments/4q2tdu/good_riddance/,self.jokes,,"I sent a reminder to a client that it was time to visit the eye doctor. He called back to inform me that he would not be coming in because, as he put it, “I have a new obstetrician.”",good riddance,1
post,4q2tcb,2qh72,jokes,false,1467025924,https://old.reddit.com/r/Jokes/comments/4q2tcb/ahahahahhaha_kia_joke_ha_yaaro/,self.jokes,,[removed],ahahahahhaha kia joke ha yaaro,0
post,4q2t30,2qh72,jokes,false,1467025795,https://old.reddit.com/r/Jokes/comments/4q2t30/did_you_know_that_the_majority_of_people_dont/,self.jokes,,[removed],Did you know that the majority of people don't know the opposite of these words?,1
post,4q2skb,2qh72,jokes,false,1467025506,https://old.reddit.com/r/Jokes/comments/4q2skb/help_ive_been_robbed/,self.jokes,,"They stole everything except my deodorant, shampoo and hand soap.

Dirty bastards ",Help! I've been robbed!,198
post,4q2s5d,2qh72,jokes,false,1467025279,https://old.reddit.com/r/Jokes/comments/4q2s5d/what_do_you_get_when_a_man_is_an_atheist_dyslexic/,self.jokes,,[deleted],"What do you get when a man is an atheist, dyslexic, and insomniac.",0
post,4q2rys,2qh72,jokes,false,1467025184,https://old.reddit.com/r/Jokes/comments/4q2rys/why_hadnt_the_law_graduate_and_the_bartender_ever/,self.jokes,,The graduate never passed the bar,Why hadn't the law graduate and the bartender ever met?,3
post,4q2rd7,2qh72,jokes,false,1467024808,https://old.reddit.com/r/Jokes/comments/4q2rd7/tommen_showed_us/,self.jokes,,[removed],Tommen showed us...,1
post,4q2r3v,2qh72,jokes,false,1467024661,https://old.reddit.com/r/Jokes/comments/4q2r3v/what_do_you_call_a_cheap_circumcision/,self.jokes,,A rip off,What do you call a cheap circumcision??,0
post,4q2qe2,2qh72,jokes,false,1467024251,https://old.reddit.com/r/Jokes/comments/4q2qe2/want_to_hear_the_funniest_joke_in_the_world/,self.jokes,,[deleted],Want to hear the funniest joke in the world?,0
post,4q2qaj,2qh72,jokes,false,1467024207,https://old.reddit.com/r/Jokes/comments/4q2qaj/wanna_here_a_joke/,self.jokes,,Britain's international trade now that they've left the EU,Wanna here a joke?,0
post,4q2ox1,2qh72,jokes,false,1467023468,https://old.reddit.com/r/Jokes/comments/4q2ox1/the_eu_now_has_1_free_gb_of_space/,self.jokes,,[removed],The EU now has 1 free 'GB' of space,1
post,4q2mqi,2qh72,jokes,false,1467022243,https://old.reddit.com/r/Jokes/comments/4q2mqi/muslims_are_like_minecraft_creepers/,self.jokes,,"If they get too close in combat, they explode 
Ps. I am Muslim ",Muslims are like minecraft creepers,0
post,4q2l5v,2qh72,jokes,false,1467021350,https://old.reddit.com/r/Jokes/comments/4q2l5v/what_is_that_italian_boy_with_two_arms_broken/,self.jokes,,He's struggling to tell his mom his need.,What is that Italian boy with two arms broken trying to do?,0
post,4q2l49,2qh72,jokes,false,1467021328,https://old.reddit.com/r/Jokes/comments/4q2l49/what_does_clint_eastwood_say_to_god_every_morning/,self.jokes,,"""Go Ahead Make My Day""",What does Clint Eastwood say to God every morning?,4
post,4q2kp9,2qh72,jokes,false,1467021093,https://old.reddit.com/r/Jokes/comments/4q2kp9/a_man_is_trying_to_get_into_a_club/,self.jokes,,[deleted],A man is trying to get into a club,0
post,4q2jgo,2qh72,jokes,false,1467020363,https://old.reddit.com/r/Jokes/comments/4q2jgo/three_fre/,self.jokes,,[removed],Three fre,1
post,4q2iie,2qh72,jokes,false,1467019838,https://old.reddit.com/r/Jokes/comments/4q2iie/roses_are_red/,self.jokes,,"Roses are red.          
         Violets are....red
          
  Tulips are red








My garden is on fire.",Roses are red,374
post,4q2hw9,2qh72,jokes,false,1467019478,https://old.reddit.com/r/Jokes/comments/4q2hw9/a_student_at_a_management_school_came_up_to_a/,self.jokes,,[removed],A student at a management school came up to a pretty girl and hugged...,1
post,4q2hpp,2qh72,jokes,false,1467019364,https://old.reddit.com/r/Jokes/comments/4q2hpp/world_war_ii_pilots_crash_on_a_deserted_island/,self.jokes,,"World War II is in full force, and a Japanese biplane and an american plane both crash after a dogfight on a deserted jungle island.

An American pilot, a German Pilot, and one Japanese pilot meet on the beach and figure they'll call a truce until they're rescued. 

""Alright you guys"" says the American. ""I'll get the fire going. You go into the forest and find anything to help set up a camp.""

The german goes off to look for food, and tells the Japanese pilot to handle the supplies. 

Time passes, and soon a roaring signal fire is going, the german pilot has returned with fruits and pig meat, but the sun is starting to go down and the Japanese soldier is nowhere to be found. 

Not wanting to be down a man in their situation, the American and the German both venture into the woods to look for him. 

They search for a long many hours and both decide to head back to camp and to continue the search tomorrow.

When they get back to their camp, the Japanese pilot jumps out from behind a rock and yells ""SUPPLIES!!!""
 ",World War II Pilots crash on a deserted island,26
post,4q2hop,2qh72,jokes,false,1467019347,https://old.reddit.com/r/Jokes/comments/4q2hop/dirty_a_man_goes_to_a_hooker/,self.jokes,,"A man goes to a $10 hooker and contracts crabs.
When he goes back to complain, the hooker laughs and says, ""What did you expect for $10? Lobsters ?""",[Dirty] A man goes to a hooker...,3
post,4q2ho9,2qh72,jokes,false,1467019342,https://old.reddit.com/r/Jokes/comments/4q2ho9/why_is_reddit_tired_of_the_broken_arms_joke/,self.jokes,,Because it appears in every mother fucking thread,Why is Reddit tired of the broken arms joke?,0
post,4q2hem,2qh72,jokes,false,1467019190,https://old.reddit.com/r/Jokes/comments/4q2hem/its_just_this_easy_to_steal_from_the_apple_store/,self.jokes,,[removed],It's just this easy to steal from the Apple Store (video),1
post,4q2hb6,2qh72,jokes,false,1467019129,https://old.reddit.com/r/Jokes/comments/4q2hb6/john_cena_develops_alzheimers/,self.jokes,,Now he's John Senile,John Cena develops Alzheimers...,0
post,4q2gxv,2qh72,jokes,false,1467018901,https://old.reddit.com/r/Jokes/comments/4q2gxv/how_do_you_spell_candy_with_two_letters/,self.jokes,,[removed],How do you spell candy with two letters?,0
post,4q2f1m,2qh72,jokes,false,1467017747,https://old.reddit.com/r/Jokes/comments/4q2f1m/til_my_housemate_doesnt_know_who_shania_twain_is/,self.jokes,,I proceeded to tell him that not knowing of her didn't impress me much...,TIL my housemate doesn't know who Shania Twain is...,0
post,4q2f01,2qh72,jokes,false,1467017722,https://old.reddit.com/r/Jokes/comments/4q2f01/a_scotsman_a_northern_irishman_and_an_englishman/,self.jokes,,[deleted],"A Scotsman, a Northern Irishman and an Englishman walk into a bar.",16
post,4q2dwn,2qh72,jokes,false,1467017061,https://old.reddit.com/r/Jokes/comments/4q2dwn/i_was_in_tesco_in_britain_this_morning/,self.jokes,,I was in tesco this morning and one of the cashiers asked the foreign couple in front of me if they wanted help packing their bags. Fuck sake love the vote was only yesterday give them a chance,I was in tesco in Britain this morning,3
post,4q2dvz,2qh72,jokes,false,1467017048,https://old.reddit.com/r/Jokes/comments/4q2dvz/dirty_joke/,self.jokes,,"An old joke I heard my dad tell my older brother years ago when I was just a little kid. Sorry if it has ever been posted before. I have never heard it anywhere else. 

So this guy gets off work and goes to a bar. He starts having a few drinks when he notices a lady across the bar watching him so he decides to go try his luck and he talks to her for a while. After a few hours and many drinks, they both decide to take a cab back to his place. 

As they arrive he struggles with the key for a moment, but as he finds success she grabs his arm and stops him. ""Wait. How you open the door will determine how the sex will turn out. If you barely open the door the sex may be too soft and will be forgettable. If you just slam the door open then the sex might be too rough and I might get hurt. How will you open the door?"" 

The guy stares at her for a few minutes before shrugging and replying ""I will probably lick the doorknob for a little while and then come in the backdoor.""",Dirty Joke,5
post,4q2du8,2qh72,jokes,false,1467017018,https://old.reddit.com/r/Jokes/comments/4q2du8/fetish/,self.jokes,,"I have a fetish for switching on air conditioning units.

It gives me vent elation.",Fetish...,3
post,4q2dtk,2qh72,jokes,false,1467017008,https://old.reddit.com/r/Jokes/comments/4q2dtk/what_happens_when_a_nectarine_is_too_tired_to/,self.jokes,,[deleted],What happens when a nectarine is too tired to take the stairs?,1
post,4q2dhn,2qh72,jokes,false,1467016819,https://old.reddit.com/r/Jokes/comments/4q2dhn/mom_dad_you_know_i_really_like_dick/,self.jokes,,[deleted],"Mom, Dad, you know I really like Dick...",0
post,4q2b95,2qh72,jokes,false,1467015535,https://old.reddit.com/r/Jokes/comments/4q2b95/little_billy_and_his_class_went_on_a_field_trip/,self.jokes,,"On their way back, the bus broke down and on top of that there was a huge storm. There was no way they could make it back that day so they decided to stay in a motel nearby for the night. The children were fed and put to bed. 

Little Billy came to Ms Marie and said he couldn't sleep and the only way he could fall asleep was to put his pinky in someone's belly button. She said, ""ok little Billy I will help you fall asleep"". So she lied beside him. After a while she had a funny feeling and  she said, ""Now there Little Billy, that ain't my belly button but something else"" and to that little Billy replied, ""Oh that's alright Ms Marie that ain't my pinky either but something else!""",Little Billy and his class went on a field trip with Ms. Marie,28
post,4q2b4v,2qh72,jokes,false,1467015462,https://old.reddit.com/r/Jokes/comments/4q2b4v/what_do_you_call_a_black_astronaut/,self.jokes,,Invisible,What do you call a black astronaut?,0
post,4q2b4a,2qh72,jokes,false,1467015451,https://old.reddit.com/r/Jokes/comments/4q2b4a/girl_with_no_arms_or_leg/,self.jokes,,"Came early, time to make a joke...So there was a girl with no arms or legs on a beach. As a man walked pass her she started crying. The man asked 'Whats the matter dear?' and the girl replied with 'I've never been hugged before.' So the man hugs her and the girl starts crying again. The man asks 'Whats wrong now?'. The girl replies with 'I've never been kissed before'. So the man kisses her and the girl starts crying yet again. So the man asks 'Whats the matter now?' The girl replies with 'I've never been fucked before.' So the man picks her up and throws her into the ocean and says 'You're fucked now.'﻿",Girl with no arms or leg,13
post,4q2b3i,2qh72,jokes,false,1467015437,https://old.reddit.com/r/Jokes/comments/4q2b3i/ice_cube_to_all_the_bregret_protest_voters/,self.jokes,,[deleted],Ice Cube to all the ''bregret'' protest voters,0
post,4q2b3b,2qh72,jokes,false,1467015432,https://old.reddit.com/r/Jokes/comments/4q2b3b/how_much_does_cersei_spend_on_fireworks/,self.jokes,,A princely sum.,How much does Cersei spend on fireworks?,0
post,4q29hi,2qh72,jokes,false,1467014535,https://old.reddit.com/r/Jokes/comments/4q29hi/bird_to_describe_trumps_penis/,self.jokes,,[deleted],Bird to describe Trump's penis.,5
post,4q29dy,2qh72,jokes,false,1467014471,https://old.reddit.com/r/Jokes/comments/4q29dy/how_many_brexiters_does_it_take_to_change_a/,self.jokes,,[deleted],How many Brexiters does it take to change a lightbulb?,0
post,4q29cz,2qh72,jokes,false,1467014455,https://old.reddit.com/r/Jokes/comments/4q29cz/a_guy_rescued_a_genie/,self.jokes,,"To return the favor, the genie offered him a wish: he could have unlimited money, or unlimited wisdom. The man chose the latter. A few days passed by, his friend came to visit him, finding him crying very fiercely and screaming the sentence: ""I should have chosen the money.""",A guy rescued a genie.,10
post,4q2999,2qh72,jokes,false,1467014400,https://old.reddit.com/r/Jokes/comments/4q2999/funny_jokes_ahahahahahahahhah/,self.jokes,,[removed],Funny Jokes AHAHAHAHAHAHAHHAH,0
post,4q297i,2qh72,jokes,false,1467014369,https://old.reddit.com/r/Jokes/comments/4q297i/how_is_batman_different_from_a_black_man/,self.jokes,,Batman can go in a store without Robin.,How is Batman different from a black man?,4
post,4q296r,2qh72,jokes,false,1467014356,https://old.reddit.com/r/Jokes/comments/4q296r/how_do_you_say_genius_sarcastically/,self.jokes,,Apple genius.,How do you say genius sarcastically?,6
post,4q293f,2qh72,jokes,false,1467014301,https://old.reddit.com/r/Jokes/comments/4q293f/feminism/,self.jokes,,[removed],Feminism.,1
post,4q28up,2qh72,jokes,false,1467014157,https://old.reddit.com/r/Jokes/comments/4q28up/how_did_our_grandparents_killed_time_when_there/,self.jokes,,"I already asked my mom, her four sisters and five brothers.",How did our grandparents killed time when there were no Smartphones and Internet?,134
post,4q27ba,2qh72,jokes,false,1467013292,https://old.reddit.com/r/Jokes/comments/4q27ba/yo_momma_so_poor/,self.jokes,,She stole macaroni from your preschool sculptures to use for dinner.,Yo momma so poor....,0
post,4q278b,2qh72,jokes,false,1467013250,https://old.reddit.com/r/Jokes/comments/4q278b/what_did_the_geologist_say_to_his_girlfriend/,self.jokes,,I am going to make the bedrock. ,What did the geologist say to his girlfriend before shagging her?,5
post,4q277r,2qh72,jokes,false,1467013240,https://old.reddit.com/r/Jokes/comments/4q277r/back_in_my_day_britain_used_to_be_part_of_the_eu/,self.jokes,,[removed],Back in my day Britain used to be part of the EU,1
post,4q26uv,2qh72,jokes,false,1467013067,https://old.reddit.com/r/Jokes/comments/4q26uv/while_getting_thrown_in_jail_my_grandmas/,self.jokes,,I guess you could say it was a cardiac arrest for battery.,"While getting thrown in jail, my grandma's pacemaker failed.",1
post,4q260f,2qh72,jokes,false,1467012617,https://old.reddit.com/r/Jokes/comments/4q260f/someone_farted_in_an_apple_store/,self.jokes,,Too bad they don't have Windows.,Someone farted in an Apple Store.,51
post,4q25z8,2qh72,jokes,false,1467012598,https://old.reddit.com/r/Jokes/comments/4q25z8/what_do_you_call_a_closet_full_of_lesbians/,self.jokes,,A liquor cabinet.,What do you call a closet full of lesbians?,3
post,4q25sn,2qh72,jokes,false,1467012506,https://old.reddit.com/r/Jokes/comments/4q25sn/a_termite_walks_into_a_bar_and_asks/,self.jokes,,"""Where is the bar tender?""",A termite walks into a bar and asks,7
post,4q25ms,2qh72,jokes,false,1467012411,https://old.reddit.com/r/Jokes/comments/4q25ms/how_many_mods_does_it_take_to_screw_in_a_light/,self.jokes,,[removed],How many mods does it take to screw in a light bulb?,10
post,4q24wf,2qh72,jokes,false,1467011996,https://old.reddit.com/r/Jokes/comments/4q24wf/what_did_one_lesbian_vampire_say_to_the_other/,self.jokes,,"""See you next month!""",What did one lesbian vampire say to the other lesbian vampire?,53
post,4q24g5,2qh72,jokes,false,1467011756,https://old.reddit.com/r/Jokes/comments/4q24g5/what_do_you_call_a_blind_dinosaur/,self.jokes,,A doyouthinkhe-saurus,What do you call a blind dinosaur?,2
post,4q24fp,2qh72,jokes,false,1467011751,https://old.reddit.com/r/Jokes/comments/4q24fp/what_is_the_difference_between_a_whale_a_shark/,self.jokes,,I don't fucking know you tell me,"What is the difference between a whale, a shark and someone from New York?",0
post,4q24ct,2qh72,jokes,false,1467011708,https://old.reddit.com/r/Jokes/comments/4q24ct/theres_some_free_space_in_the_eu_now1_gb_to_be/,self.jokes,,[removed],"There's some free space in the EU now....1 GB, to be precise...😊",0
post,4q22de,2qh72,jokes,false,1467010678,https://old.reddit.com/r/Jokes/comments/4q22de/how_hot_is_it/,self.jokes,,[removed],How hot is it?,1
post,4q211p,2qh72,jokes,false,1467009952,https://old.reddit.com/r/Jokes/comments/4q211p/how_do_you_piss_off_someone_on_reddit/,self.jokes,,[removed],How do you piss off someone on reddit?,1
post,4q2109,2qh72,jokes,false,1467009923,https://old.reddit.com/r/Jokes/comments/4q2109/three_large_girls_walk_into_a_bar/,self.jokes,,"They sit down at the bar and try to order a drink. The bartender clearly doesn't understand their heavy accents so a man comes over to try and help. The man says, ""excuse me, but are you ladies from Scotland?"" 

They say, ""No! Wales, Wales!""

""Oh my apologies! Are you whales from Scotland?""",Three large girls walk into a bar...,25
post,4q1zn6,2qh72,jokes,false,1467009223,https://old.reddit.com/r/Jokes/comments/4q1zn6/i_discovered_recently_that_i_can_cut_wood_just_by/,self.jokes,,It's true I saw it with my eyes,I discovered recently that I can cut wood just by looking at it,107
post,4q1z4n,2qh72,jokes,false,1467008959,https://old.reddit.com/r/Jokes/comments/4q1z4n/what_do_you_get_when_you_combine_reddit_with_dry/,self.jokes,,Circle jerky.,What do you get when you combine Reddit with dry humor?,2
post,4q1xi7,2qh72,jokes,false,1467008070,https://old.reddit.com/r/Jokes/comments/4q1xi7/my_iguana/,self.jokes,,My Iguana has been having trouble getting enough blood into his weenus; he has areptile dysfunction.,My Iguana,2
post,4q1w4y,2qh72,jokes,false,1467007370,https://old.reddit.com/r/Jokes/comments/4q1w4y/this_is_the_latest_trend_for_timepass_follow_this/,self.jokes,,[removed],This is the latest trend for TIMEPASS !!! Follow this popular &amp; clean Telegram channel.,1
post,4q1vz9,2qh72,jokes,false,1467007289,https://old.reddit.com/r/Jokes/comments/4q1vz9/a_man_walks_into_a_library_and_says_to_the/,self.jokes,,"The librarian looks on her computer and says, ""I don't know if it's in yet.""
""Yeah that's the one""","A man walks into a library and says to the librarian, ""do you have that book for men with small penises?""",155
post,4q1vyw,2qh72,jokes,false,1467007283,https://old.reddit.com/r/Jokes/comments/4q1vyw/why_was_six_afraid_of_seven/,self.jokes,,Because seven was a registered child molester.,Why was six afraid of seven?,10
post,4q1vwd,2qh72,jokes,false,1467007244,https://old.reddit.com/r/Jokes/comments/4q1vwd/what_do_cannibals_call_plane_crash_victims/,self.jokes,,[deleted],What do cannibals call plane crash victims?,0
post,4q1vhi,2qh72,jokes,false,1467007034,https://old.reddit.com/r/Jokes/comments/4q1vhi/what_do_you_call_a_nice_canadian_meal_on_a/,self.jokes,,Poutina.,What do you call a nice Canadian meal on a colorful roof?,0
post,4q1vbg,2qh72,jokes,false,1467006951,https://old.reddit.com/r/Jokes/comments/4q1vbg/why_did_the_firemen_go_to_the_classroom/,self.jokes,,It was a heated debate.,Why did the firemen go to the classroom?,1
post,4q1v6h,2qh72,jokes,false,1467006878,https://old.reddit.com/r/Jokes/comments/4q1v6h/knock_knock/,self.jokes,,"""who's there?"" 

""Europe""

""Europe who?""

""No, you're a poo""",Knock knock,0
post,4q1uy2,2qh72,jokes,false,1467006754,https://old.reddit.com/r/Jokes/comments/4q1uy2/build_a_man_a_fire_and_you_warm_him_for_a_day/,self.jokes,,Light a man on fire and you warm him for the rest of his life.,Build a man a fire and you warm him for a day.,81
post,4q1uss,2qh72,jokes,false,1467006683,https://old.reddit.com/r/Jokes/comments/4q1uss/a_koala_was_sitting_in_a_tree_smoking_a_joint/,self.jokes,,[deleted],A koala was sitting in a tree smoking a joint...,0
post,4q1uij,2qh72,jokes,false,1467006537,https://old.reddit.com/r/Jokes/comments/4q1uij/if_i_had_a_dollar_for_every_joke_ive_recycled/,self.jokes,,I would have a lot since this is a popular style of joke,If I had a dollar for every joke I've recycled,2
post,4q1uc9,2qh72,jokes,false,1467006445,https://old.reddit.com/r/Jokes/comments/4q1uc9/what_do_teenage_terrorists_drink/,self.jokes,,Smirnoff ISIS,What do teenage terrorists drink?,1
post,4q1u5o,2qh72,jokes,false,1467006340,https://old.reddit.com/r/Jokes/comments/4q1u5o/a_trip_to_wales/,self.jokes,,"A couple are driving through Wales late one night and they pass through Llanfairpwllgwyngyllgogerychwyrndrobwilllantysiliogogogoch. With nothing much else to do , they start arguing over the pronunciation. Eventually they decide to stop somewhere and ask a local. They pull up somewhere and go inside, and ask the staff member ""excuse me, could you pronounce the name of this place, really slowly?""
The kid behind the counter gives them a confused look, and says ""burr-gurr kiiiiing""",A trip to Wales.,77
post,4q1sw9,2qh72,jokes,false,1467005711,https://old.reddit.com/r/Jokes/comments/4q1sw9/how_does_a_welshman_find_sheep_in_tall_grass/,self.jokes,,Irresistible.,How does a Welshman find sheep in tall grass?,9
post,4q1sc4,2qh72,jokes,false,1467005465,https://old.reddit.com/r/Jokes/comments/4q1sc4/a_woman_is_going_into_labor/,self.jokes,,"... so the husband and wife quickly head to the hospital.  After they arrive the doctor comes into the room and says to the couple, ""We have developed a new experimental treatment where we can hook you up to a machine and transfer some of the pain from labor to the father.  I warn you though that even 10% transference will be the most pain he has ever felt before in his life.""  The husband, not wanting his wife to suffer, said okay to the treatment.  So the doctor hooks the woman up to the machine and turns it on to 5% just to start.  After a few minutes of waiting he asks the husband if he's okay to increase the percentage and he says yes.  The doctor continues to crank it up to 10% and again asks the husband if he's okay and again the husband says that he's fine. The doctor, a little confused now, turns the machine up higher to 50%.  The husband still says that he's fine and the wife seems to be feeling much less pain. The doctor, completely bewildered now, cranks the machine all the way up to 100% and the baby is delivered relatively pain free and the couple go home.

When they get home the mail man is dead on the porch.",A Woman Is Going Into Labor,0
post,4q1s7x,2qh72,jokes,false,1467005411,https://old.reddit.com/r/Jokes/comments/4q1s7x/why_are_gametes_best_suited_to_advertising_careers/,self.jokes,,Because sex cells.,Why are gametes best suited to advertising careers?,13
post,4q1rse,2qh72,jokes,false,1467005216,https://old.reddit.com/r/Jokes/comments/4q1rse/has_anyone_else_realized/,self.jokes,,that sierra mist and mountain dew are technically the same thing,Has anyone else realized...,0
post,4q1qtb,2qh72,jokes,false,1467004771,https://old.reddit.com/r/Jokes/comments/4q1qtb/two_american_soldiers_have_taken_cover_in_a/,self.jokes,,"The enemy fire power is fierce, and they are unable to advance or retreat.  Shells are zinging past them like wasps, and errant ricochets unnerve them.    Mortar shells explode all around and the two men are sweating lest a shell might land atop of them.  As the evening wears on and nerves become frazzled in the stifling heat, one of the men confides that he has to go to the bathroom really bad.  ""Number  1 or Number 2?"" his friend asks.  ""Number 2.""  He says.  ""Well you can't do your business in here.  There is no telling how long we'll be trapped in this foxhole before reinforcements arrive to liberate us.  So you'll just have to hold it.""

Nighttime falls, but the shelling does not let up.  With daylight the two men peer outside to discover it would be another long day of hunkering down.   As the minutes build into hours the one soldier finally blurts out, ""Joe, I just can't hold it any longer.  I've gotta go to the bathroom.""  Joe looks over at his companion who is ashen faced, and visibly sweating:  ""Well Slim, it appears that you have two choices.  Take a crap in here and I shoot you, or go and do it out there and the Germans shoot you.  Which will it be?""

""I've been considering that,"" says Slim.  ""Do you see that foxhole over  yonder?""  and he points it out.  ""I saw a mortar shell land atop of it yesterday and there's been no activity since, so I can safely say the fellas inside won't complain if I use it as a latrine.  If you'll cover me, I think I can make it over , do my business, signal you, and then come back under your cover fire.""

Joe agrees, and Slim makes a successful dash for the neighboring foxhole while he lays down the cover fire.  ""Damn if the lucky fool didn't make it,"" Joe swore.  Half an hour passed as Joe waited for the signal from Slim.  No Slim.  An hour passed.  Still no Slim.  Two hours.  Then Three hours.  No Slim.  Nightfall arrived and still no signal came from the other foxhole.  ""I guess Ol' Slim must have caught a bullet after all.""  He  said remorsefully, and turned in for the night.

Come daylight, Joe's eyes were on the neighboring foxhole intently hoping for a signal from his friend.  It never came.  That day too passed as uneventfully as the one before it, and Joe was convinced Slim was dead.   But come the next morning, Joe was amazed to see Slim signaling at him from the neighboring foxhole.  Joe signaled back, and laid down a cover fire as Slim made his mad dash back.  Diving inside just as a cavalcade of enemy bullets smashed into the sandbags.

""What the hell took you so long over there?""  Joe asked.

""You wouldn't believe me if I told you,"" said Slim.

""Try me.""  Says Joe.

""Well pard, when I dove into that foxhole.  I landed right on top of one of them Red Cross nurses.  Her name was Sally, and she must be around nineteen years old, and her with the best figure I've seen on a woman since this war started.""

""Damn your luck,""  says Joe.  ""What'd you do.""

""What do you think?""  Slim answered.  ""I was a man, she was a woman.    We have been making sweet. sweet love from that moment on.""

""You have been making love this entire time?""  Joe asks.

""Damn straight.""  Slim says.   

""Hot damn!""  Joe stutters.  ""Do you suppose she'll be willing to give me a roll in the hay if I was to make a call over to that foxhole myself.""

""She's not a woman to turn a man down, that's for sure.""  Assures Slim.

""Oh boy.  Oh boy.""  Says Joe as sheds his heavy backpack.  ""You say she has a shapely figure.  How is she for looks?""

""You know what pard,"" Slim answers.  ""I couldn't rightly say.  That damn mortar had taken her head clean off.""
",Two American soldiers have taken cover in a foxhole during an offensive in France during ww2.,4
post,4q1qrf,2qh72,jokes,false,1467004747,https://old.reddit.com/r/Jokes/comments/4q1qrf/girl_making_sandwich/,self.jokes,,[removed],Girl making sandwich,1
post,4q1pui,2qh72,jokes,false,1467004327,https://old.reddit.com/r/Jokes/comments/4q1pui/a_few_years_ago_i_was_at_the_pub_sitting_at_the/,self.jokes,,"Being new to the area and friendly, I say ""Oh! Are you two ladies from England?""

The one closest to me gets a look of disgust and with a super bitchy tone says ""Actually, it's Wales"".

So I reply ""Oh, I'm sorry. Are you two whales from England?""",A few years ago I was at the pub. Sitting at the end of the bar were two large middle-aged women speaking in what I thought were thick English accents.,4
post,4q1ppc,2qh72,jokes,false,1467004264,https://old.reddit.com/r/Jokes/comments/4q1ppc/john_and_peter/,self.jokes,,"John: Dude my girlfriend is pregnant, but I use a condom every time.

Peter: Come here my dear friend and I will explain it to you

John: Ok.

Peter: A man went into the jungle with an umbrella. He saw a tiger coming right at him. He touched the button of his umbrella and the tiger died. 

John: Haha!But that's impossible. Maybe someone else shot the tiger.

Peter: Exactly..
",John and Peter,24
post,4q1oi5,2qh72,jokes,false,1467003748,https://old.reddit.com/r/Jokes/comments/4q1oi5/what_is_lionel_messis_favorite_soft_drink/,self.jokes,,"Si, era Missed",What is Lionel Messi's favorite soft drink?,4
post,4q1oau,2qh72,jokes,false,1467003651,https://old.reddit.com/r/Jokes/comments/4q1oau/what_did_the_communist_pig_call_his_writings/,self.jokes,,[deleted],what did the communist pig call his writings?,6
post,4q1o0u,2qh72,jokes,false,1467003516,https://old.reddit.com/r/Jokes/comments/4q1o0u/why_are_crabs_always_so_tired/,self.jokes,,It's because they only sleep in snatches.,Why are crabs always so tired?,1
post,4q1mvq,2qh72,jokes,false,1467002961,https://old.reddit.com/r/Jokes/comments/4q1mvq/teacher_asks_johnny_whats_wrong/,self.jokes,,"Johnny :- Our house is very small. Me, my mum and my dad sleep on the same bed. Every night my dad asks, 'Johnny, are you asleep?'

I say No &amp; he slaps my face &amp; gives me a Black eye

Teacher:- Tonight, when your dad asks again, keep dead quiet &amp; don't answer.

The following morning Johnny comes back with a severe black eye again.

Teacher:- My goodness why the black eye again? Johnny:- Dad asked me if I was asleep. I shut up &amp; kept dead still. Then my mum and dad started moving at the same time. Mum was breathing erratically, kicking her legs up frantically &amp; squealing like a hyena on the bed. Then my dad asked my mum, ""Are you coming?"" Mum said, ""Yes I'm coming, are you coming too?"" Dad answered:- Yes.

Well, they don't usually go anywhere without me so I said, ""wait for me, I'm coming too"".
","Teacher asks Johnny, ""What's Wrong?""",165
post,4q1l2n,2qh72,jokes,false,1467002164,https://old.reddit.com/r/Jokes/comments/4q1l2n/where_was_mercy_during_the_holocaust/,self.jokes,,[removed],Where was Mercy during the Holocaust?,1
post,4q1kt5,2qh72,jokes,false,1467002052,https://old.reddit.com/r/Jokes/comments/4q1kt5/a_condom_doesnt_guarantee_safe_sex/,self.jokes,,My friend was wearing one when he was shot by the woman's husband.,A condom doesn't guarantee safe sex.,4
post,4q1kc9,2qh72,jokes,false,1467001843,https://old.reddit.com/r/Jokes/comments/4q1kc9/computer_nerd_dirty_talk/,self.jokes,,I'm going to stick my D: disk into your V: drive.,Computer nerd dirty talk,0
post,4q1k55,2qh72,jokes,false,1467001773,https://old.reddit.com/r/Jokes/comments/4q1k55/my_girlfriend_says_she_prefers_a_dildo_over_me/,self.jokes,,I never saw it coming,My girlfriend says she prefers a dildo over me.,10
post,4q1jne,2qh72,jokes,false,1467001573,https://old.reddit.com/r/Jokes/comments/4q1jne/a_teacher_comes_to_a_students_house_for_a_parent/,self.jokes,,"A teacher comes over to a student's house for a parent teacher meeting. The mom is making turkey in the kitchen and the dad is shaving for the occasion. The teacher rings the doorbell and the student answers and allows the teacher to come in. The teacher asks, ""What are your parents doing?"" The student goes to check in on his mom first. While cutting the turkey the mom cuts a finger and yells ""**FUCK!**"" Then the student goes to the bathroom to see how his dad is doing. The Dad cuts himself while shaving and yells ""**SHIT!**"" The student then comes back down and tells the teacher, ""My mom is fucking a turkey in the kitchen and my dad is shitting himself in the bathroom.""",A teacher comes to a student's house for a parent teacher meeting,0
post,4q1iqi,2qh72,jokes,false,1467001126,https://old.reddit.com/r/Jokes/comments/4q1iqi/how_many_suh_goods_does_it_take_to_screw_in_a/,self.jokes,,none its already lit sam hahahah ssoooohh,How many 'suh goods' does it take to screw in a light bulb?,0
post,4q1hjy,2qh72,jokes,false,1467000601,https://old.reddit.com/r/Jokes/comments/4q1hjy/why_did_the_operation_barbarossa_fail/,self.jokes,,The supreme commander didn't have the balls required.,Why did the operation Barbarossa fail?,0
post,4q1h5s,2qh72,jokes,false,1467000413,https://old.reddit.com/r/Jokes/comments/4q1h5s/did_you_hear_about_the_man_who_was_arrested_for/,self.jokes,,He was suspected of Fowl Play,Did you hear about the man who was arrested for molesting a duck?,20
post,4q1gex,2qh72,jokes,false,1467000109,https://old.reddit.com/r/Jokes/comments/4q1gex/tonight_on_my_strange_addition/,self.jokes,,Man addicted to brake fluid claims he can stop at any time,Tonight on My Strange Addition,0
post,4q1fwl,2qh72,jokes,false,1466999899,https://old.reddit.com/r/Jokes/comments/4q1fwl/it_is_said_that_wearing_tshirts_make_you_feel/,self.jokes,,I've been wearing a dozen of them but it's still hot like hell. Damn.,It is said that wearing T-shirts make you feel cooler in Summer,10
post,4q1fmu,2qh72,jokes,false,1466999788,https://old.reddit.com/r/Jokes/comments/4q1fmu/did_anyone_see_got_tonight_spoilers/,self.jokes,,Tommen took King's Landing much too seriously,Did anyone see GOT tonight? (spoilers!!!),1
post,4q1f7l,2qh72,jokes,false,1466999610,https://old.reddit.com/r/Jokes/comments/4q1f7l/what_did_ser_gayme_lannister_name_his_dong/,self.jokes,,[deleted],What did Ser Gayme Lannister name his dong?,1
post,4q1eya,2qh72,jokes,false,1466999514,https://old.reddit.com/r/Jokes/comments/4q1eya/there_is_a_man_with_a_friend_who_is_a_ninja/,self.jokes,,"The man asks, ""Ninja, can you help me out with this lightbulb?""


The ninja replies ""Shur-i-ken!""",There is a man with a friend who is a ninja....,4
post,4q1etg,2qh72,jokes,false,1466999463,https://old.reddit.com/r/Jokes/comments/4q1etg/in_the_future_a_group_of_scientists_invent_a_very/,self.jokes,,[deleted],"In the future, a group of scientists invent a very powerful computer",2
post,4q1e8j,2qh72,jokes,false,1466999205,https://old.reddit.com/r/Jokes/comments/4q1e8j/little_april_was_not_the_best_student_in_sunday/,self.jokes,,"Little April was not the best student in Sunday school. Usually she slept through the class. One day the teacher called on her while she was napping, ""Tell me, April, who created the universe?"" When April didn't stir, little Johnny, a boy seated in the chair behind her, took a pin and jabbed her in the rear. ""GOD ALMIGHTY!"" shouted April and the teacher said, ""Very good"" and April fell back asleep. A while later the teacher asked April, ""Who is our Lord and Saviour,"" But, April didn't even stir from her slumber. Once again, Johnny came to the rescue and stuck her again. ""JESUS CHRIST!"" shouted April and the teacher said, ""very good,"" and April fell back to sleep. Then the teacher asked April a third question. ""What did Eve say to Adam after she had her twenty-third child?"" And again, Johnny jabbed her with the pin. This time April jumped up and shouted, ""IF YOU STICK THAT F*****G THING IN ME ONE MORE TIME, I'LL BREAK IT IN HALF AND STICK IT UP YOUR ARSE!"" The Teacher fainted.",Little April was not the best student in Sunday school,63
post,4q1e1f,2qh72,jokes,false,1466999126,https://old.reddit.com/r/Jokes/comments/4q1e1f/what_happens_when_you_put_nutella_on_salmon/,self.jokes,,[deleted],What happens when you put nutella on salmon?,0
post,4q1dr7,2qh72,jokes,false,1466999005,https://old.reddit.com/r/Jokes/comments/4q1dr7/how_do_you_know_if_your_car_is_gay/,self.jokes,,[deleted],How do you know if your car is gay?,0
post,4q1dez,2qh72,jokes,false,1466998864,https://old.reddit.com/r/Jokes/comments/4q1dez/an_girl_cooks_for_her_exboyfriend/,self.jokes,,"The girl cooks a dish for her ex-boyfriend. He takes a bite.

The girl asks, ""What does it taste like""

The boy says, ""It tastes like your personality.""",An girl cooks for her ex-boyfriend...,0
post,4q1ckr,2qh72,jokes,false,1466998515,https://old.reddit.com/r/Jokes/comments/4q1ckr/so_a_newly_wed_couple_is_about_to_have_their/,self.jokes,,[deleted],So a newly wed couple is about to have their first night...,0
post,4q1c0b,2qh72,jokes,false,1466998289,https://old.reddit.com/r/Jokes/comments/4q1c0b/in_the_year_2060/,self.jokes,,"In the year 2060, owning guns has been outlawed. Men and women clothed in black armor approach a small cottage. Inside the cottage is a man with a grey beard and a glass of scotch. One of the soldiers kicks down the old wooden door and proclaims, ""We're here for your arms!"" The Old man sits quietly, picks up the glass of scotch, and takes a swig. ""You can't have my arms, I need them to eat and drink.""",In the year 2060,0
post,4q1bwh,2qh72,jokes,false,1466998242,https://old.reddit.com/r/Jokes/comments/4q1bwh/why_did_lionel_messi_cross_the_road/,self.jokes,,to retrieve his penalty kick ,Why did Lionel Messi cross the road?,1
post,4q1b14,2qh72,jokes,false,1466997886,https://old.reddit.com/r/Jokes/comments/4q1b14/america_and_britain_are_in_the_having_a/,self.jokes,,[removed],America and Britain are in the having a competition on who can fuck themselves up the most.,0
post,4q19zq,2qh72,jokes,false,1466997471,https://old.reddit.com/r/Jokes/comments/4q19zq/whats_the_difference_between_a_catholic_priest/,self.jokes,,A pimple doesn't come on a boys face until he's 13,What's the difference between a Catholic priest and a pimple?,33
post,4q19kf,2qh72,jokes,false,1466997303,https://old.reddit.com/r/Jokes/comments/4q19kf/on_a_scale_of_gorilla_to_alligator_how_shitty_of/,self.jokes,,[removed],On a scale of gorilla to alligator... How shitty of a parent are you?,1
post,4q18zk,2qh72,jokes,false,1466997061,https://old.reddit.com/r/Jokes/comments/4q18zk/how_do_you_lose_a_football_championship_penalty/,self.jokes,,You Messi-up,How do you lose a Football championship penalty shootout?,0
post,4q18r5,2qh72,jokes,false,1466996981,https://old.reddit.com/r/Jokes/comments/4q18r5/did_you_hear_how_argentina_lost_the_game/,self.jokes,,heard it was pretty Messi,Did you hear how Argentina lost the game?,2
post,4q17dl,2qh72,jokes,false,1466996462,https://old.reddit.com/r/Jokes/comments/4q17dl/so_a_mexican_sneaks_across_the_border_into_america/,self.jokes,,"And the border patrol officer says ""Oh no not again""",So a Mexican sneaks across the border into America,0
post,4q15sh,2qh72,jokes,false,1466995853,https://old.reddit.com/r/Jokes/comments/4q15sh/game_of_thrones_season_6_finale_spoiler_what/,self.jokes,,[removed],[Game of Thrones Season 6 finale spoiler] What would you call the aftermath of that one character's suicide?,0
post,4q15e7,2qh72,jokes,false,1466995698,https://old.reddit.com/r/Jokes/comments/4q15e7/so_a_man_goes_on_a_date/,self.jokes,,"And says, ""I hope you don't mind I brought my mother along."" to his date.
She says, ""Ummm...it's ok I guess, where is she?""
He places an urn on table, and says:
""Mom this is Laura, Laura this is my mom, Cathy.""",So a man goes on a date...,0
post,4q158c,2qh72,jokes,false,1466995635,https://old.reddit.com/r/Jokes/comments/4q158c/i_dont_like_male_pornstars/,self.jokes,,They always are fucking assholes,I don't like male pornstars,1
post,4q14uk,2qh72,jokes,false,1466995486,https://old.reddit.com/r/Jokes/comments/4q14uk/when_im_stressed_i_go_to_the_gym/,self.jokes,,Cause then I could workout my problems,"When I'm stressed, I go to the gym",0
post,4q13zy,2qh72,jokes,false,1466995170,https://old.reddit.com/r/Jokes/comments/4q13zy/how_do_you_know_when_a_woman_is_about_to_say_some/,self.jokes,,"She starts her sentance with ""A man once told me""",How do you know when a woman is about to say some thing intelligent?,4
post,4q138b,2qh72,jokes,false,1466994889,https://old.reddit.com/r/Jokes/comments/4q138b/hilary_clinton_might_become_the_first_f_president/,self.jokes,,[deleted],Hilary Clinton might become the first F president...,0
post,4q130q,2qh72,jokes,false,1466994803,https://old.reddit.com/r/Jokes/comments/4q130q/so_i_guess_the_eu/,self.jokes,,I guess the EU has 1 GB of free space now ,So I guess the EU,4
post,4q12wt,2qh72,jokes,false,1466994761,https://old.reddit.com/r/Jokes/comments/4q12wt/america_and_britain_are_having_a_competition/,self.jokes,,"To see who can fuck themselves up the most. 

Britain is currently winning, but the USA has a Trump card.",America and Britain are having a competition,0
post,4q12up,2qh72,jokes,false,1466994741,https://old.reddit.com/r/Jokes/comments/4q12up/what_field_of_study_did_the_pirate_accountant_get/,self.jokes,,[deleted],What field of study did the pirate accountant get into?,0
post,4q12mx,2qh72,jokes,false,1466994655,https://old.reddit.com/r/Jokes/comments/4q12mx/what_do_you_call_a_blueeyed_blonde_that_doesnt/,self.jokes,,A vegetaryan,What do you call a blue-eyed blonde that doesn't eat meat?,30
post,4q124y,2qh72,jokes,false,1466994465,https://old.reddit.com/r/Jokes/comments/4q124y/whats_the_best_way_to_sum_up_the_90s/,self.jokes,,90+91+92+93+94+95+96+97+98+99=945,What's the best way to sum up the 90's?,132
post,4q11ep,2qh72,jokes,false,1466994192,https://old.reddit.com/r/Jokes/comments/4q11ep/cah_online/,self.jokes,,[removed],CAH Online,1
post,4q119a,2qh72,jokes,false,1466994138,https://old.reddit.com/r/Jokes/comments/4q119a/spoiler_if_you_watched_game_of_thrones/,self.jokes,,[deleted],[Spoiler] If you watched Game of Thrones,1
post,4q0zye,2qh72,jokes,false,1466993628,https://old.reddit.com/r/Jokes/comments/4q0zye/what_drugs_do_cows_take/,self.jokes,,Cow-caine,What drugs do cows take?,0
post,4q0zv0,2qh72,jokes,false,1466993587,https://old.reddit.com/r/Jokes/comments/4q0zv0/fun_facts/,self.jokes,,"The reason that their are only 49 contestants in the Miss America Contest is because nobody wants to wear a banner that says ""IDAHO""

My mind is like a bear trap. Rusty and illegal in 37 states.

My neighbour knocked on my door at 2 AM! Can you believe it? He's lucky I was up playing with my Heavy Metal band!

Every day, you beat your previous record of consecutive days alive.

Fire fighting is like sex - The most important things are Size, equipment and technique.

Politicians and diapers have a lot in common. They both should be changed frequently, and for the same reason. ",Fun Facts,15
post,4q0xy8,2qh72,jokes,false,1466992787,https://old.reddit.com/r/Jokes/comments/4q0xy8/after_years_in_the_military/,self.jokes,,"After years in the Military, the soldier survived mustard gas and pepper spray and was proud to finally be able to call himself a seasoned veteran.",After years in the Military,89
post,4q0xsf,2qh72,jokes,false,1466992720,https://old.reddit.com/r/Jokes/comments/4q0xsf/ive_got_99_problems/,self.jokes,,[deleted],I've got 99 problems...,1
post,4q0xhg,2qh72,jokes,false,1466992597,https://old.reddit.com/r/Jokes/comments/4q0xhg/my_vacation/,self.jokes,,[deleted],my vacation,1
post,4q0xad,2qh72,jokes,false,1466992506,https://old.reddit.com/r/Jokes/comments/4q0xad/best_exercise_to_lose_a_few_pounds/,self.jokes,,"So my friend who is a fitness instructor just came up with a new exercise to lose pounds in just a matter of days. He calls it the ""Brexit"".",Best exercise to lose a few pounds...,29
post,4q0wt5,2qh72,jokes,false,1466992298,https://old.reddit.com/r/Jokes/comments/4q0wt5/three_econometricians_went_out_hunting_and_came/,self.jokes,,"The first econometrician fired, but missed by one meter to the left. The second econometrician fire, but missed by one meter to the right. The third econometrician didn't fire, but shouted in triumph, ""We got it! We got it!""",Three econometricians went out hunting and came across a large deer.,9
post,4q0wj5,2qh72,jokes,false,1466992180,https://old.reddit.com/r/Jokes/comments/4q0wj5/a_man_comes_home_from_work_and_says_to_his_wife/,self.jokes,,"""What do you think? Is that something you could get behind?""","A man comes home from work and says to his wife, ”Honey, I'm thinking about ordering a strap-on dildo from Amazon...""",5
post,4q0wfg,2qh72,jokes,false,1466992137,https://old.reddit.com/r/Jokes/comments/4q0wfg/lol/,self.jokes,,[removed],LOL,1
post,4q0w2x,2qh72,jokes,false,1466991984,https://old.reddit.com/r/Jokes/comments/4q0w2x/why_cant_america_play_chess/,self.jokes,,They are missing 2 towers,Why can't America play chess?,34
post,4q0vy2,2qh72,jokes,false,1466991922,https://old.reddit.com/r/Jokes/comments/4q0vy2/what_did_samuel_l_jackson_say_when_he_saw_a_guy/,self.jokes,,[deleted],What did Samuel L. Jackson say when he saw a guy being eaten by a velociraptor?,0
post,4q0vn2,2qh72,jokes,false,1466991795,https://old.reddit.com/r/Jokes/comments/4q0vn2/setting_up_a_sexual_innuendo_club/,self.jokes,,"Let me know if you can come! It will be a bit hard to set up, but to give it to you straight, I'm sure it will leave you satisfied and smiling!
Wood you mind telling your friends? Feel free to accept, since you can always just pull out!",Setting up a Sexual Innuendo club,0
post,4q0vjh,2qh72,jokes,false,1466991755,https://old.reddit.com/r/Jokes/comments/4q0vjh/what_disease_does_jar_jar_binks_get_after_he_is/,self.jokes,,[deleted],What disease does Jar Jar Binks get after he is exposed to asbestos?,1
post,4q0v2t,2qh72,jokes,false,1466991566,https://old.reddit.com/r/Jokes/comments/4q0v2t/my_friend_recently_died_from_aids_that_he/,self.jokes,,At least he died doing what he loved.,My friend recently died from AIDS that he contracted from his partner,0
post,4q0umt,2qh72,jokes,false,1466991386,https://old.reddit.com/r/Jokes/comments/4q0umt/a_guy_walks_up_to_a_girl_in_the_bar_with_his_fist/,self.jokes,,"The girl says........The empire state building.

The guy says..........That's close enough.",A guy walks up to a girl in the bar with his fist closed and says........I will go down on you if you can guess what I have in my hand.,45
post,4q0ubg,2qh72,jokes,false,1466991265,https://old.reddit.com/r/Jokes/comments/4q0ubg/have_you_ever_been_to_a_native_american_orgy/,self.jokes,,It's fucking intense man!,Have you ever been to a Native American orgy?,0
post,4q0tw9,2qh72,jokes,false,1466991099,https://old.reddit.com/r/Jokes/comments/4q0tw9/how_do_you_say_virgin_in_dutch/,self.jokes,,Goodentight,"How do you say ""virgin"" in Dutch?",2
post,4q0ror,2qh72,jokes,false,1466990184,https://old.reddit.com/r/Jokes/comments/4q0ror/there_wasnt_much_time_left_the_man_had_to_act/,self.jokes,,[deleted],There wasn't much time left - the man had to act quickly.,5
post,4q0r6j,2qh72,jokes,false,1466989962,https://old.reddit.com/r/Jokes/comments/4q0r6j/hey_dad_did_you_get_a_haircut/,self.jokes,,"No son, I got all of 'em cut","Hey dad, did you get a haircut?",0
post,4q0qe0,2qh72,jokes,false,1466989663,https://old.reddit.com/r/Jokes/comments/4q0qe0/did_you_know_that_the_majority_of_people_dont/,self.jokes,,[deleted],Did you know that the majority of people don't know the opposite of these words?,10776
post,4q0pse,2qh72,jokes,false,1466989417,https://old.reddit.com/r/Jokes/comments/4q0pse/why_did_lucy_fall_off_the_swing/,self.jokes,,"Jimmy pushed her...

Which is a shame because she was getting used to swinging without arms.",Why did Lucy fall off the swing?,0
post,4q0otj,2qh72,jokes,false,1466989016,https://old.reddit.com/r/Jokes/comments/4q0otj/my_left_butt_cheek_was_hurting_pretty_bad_earlier/,self.jokes,,that I didn't want it half-assed.,"My left butt cheek was hurting pretty bad earlier, so I asked my girlfriend to massage it for me. I told her...",7
post,4q0ogu,2qh72,jokes,false,1466988866,https://old.reddit.com/r/Jokes/comments/4q0ogu/whats_the_difference_between_the_mailman_and_the/,self.jokes,,The mailman doesn't come on Sunday.,What's the difference between the mailman and the priest?,0
post,4q0o27,2qh72,jokes,false,1466988683,https://old.reddit.com/r/Jokes/comments/4q0o27/making_english_the_language_of_the_eu/,self.jokes,,"The European Commission have just announced an agreement whereby English will be the official language of the EU rather than German, which was the other possibility. As part of the negotiations, Her Majesty's govt. conceded that English spelling had some room for improvement and has accepted a 5 year phase in plan that would be known as ""EuroEnglish"".

In the first year, ""s"" will replace the soft ""c"".. Sertainly, this will make the sivil servants jump with joy. The hard ""c"" will be dropped in favor of the ""k"". This should klear up konfusion and keyboards kan have 1 less letter.

There will be growing publik enthusiasm in the sekond year, when the troublesome  ""ph"" will be replaced with the ""f"". This will make words like ""fotograf"" 20% shorter.

In the 3rd year, publik akseptanse of the new spelling kan be expekted to reach the stage where more komplikated changes are possible. Governments will enkorage the removal of double letters, which have always ben a deterent to akurate speling. Also, al wil agre  that the horible mes of the silent ""e""'s in the language is disgraceful, and they should go away.

By the 4th yar, peopl wil be reseptiv to steps such as replasing ""th"" with ""z"" and ""w"" with ""v"".

During ze fifz year, ze unesesary ""o"" kan be dropd from vords kontaining ""ou"" and similar changes vud of kors be aplid to ozer kombinations of leters.

After zis fifz yer, ve vil hav a reli sensibl riten styl. Zer vil be no mor trubls or difikultis and evrivun vil find it ezi tu understand ech ozer.

ZEN ZE DREM VIL FINALI KUM TRU!! And zen ve vil take over ze vorld!!!
",Making English the language of the EU,10
post,4q0nvj,2qh72,jokes,false,1466988603,https://old.reddit.com/r/Jokes/comments/4q0nvj/a_doctor_tries_to_make_some_money_off_of_an/,self.jokes,,"An unemployed engineer who was tired of being jobless opens his own medical clinic. ""A cure for your ailment guaranteed at $500; we'll play you $1,000 if we fail.""
A doctor thinks this is a good opportunity to earn $1,000, and goes to the clinic.

Doctor: ""I have lost my sense of taste.""

Engineer: ""Nurse, please bring the medicine from box 22 and put 3 drops in the patient's mouth.""

Doctor: ""This is gasoline!""

Engineer: ""Congratulations! You've got your taste back. That will be $500.""

The doctor gets annoyed and goes back to a couple days to hopefully recover his money.

Doctor: ""I have lost my memory, I can't remember anything!""

Engineer: ""Nurse please bring the medicine from box 22 and put 3 drops in the patients mouth.""

Doctor: ""But that's gasoline!""

Engineer: ""Congratulations! You've got your memory back. That will me $500.""

The doctor leaves angrily, but returns several days later more determined than every to make is money back. 

Doctor: ""I've lost my eyesight.""

Engineer: ""Well I don't have any cure for this. Take this $1,000,"" passing the doctor only $500.

Doctor: ""But this is only $500!""

Engineer: ""Congratulations! You've got your eyesight back. That will me $500.""",A Doctor tries to make some money off of an engineer,71
post,4q0nr6,2qh72,jokes,false,1466988551,https://old.reddit.com/r/Jokes/comments/4q0nr6/what_did_the_sperm_say_to_the_egg/,self.jokes,,Nice to meet you. Wanna make a baby?,What did the sperm say to the egg?,0
post,4q0noj,2qh72,jokes,false,1466988515,https://old.reddit.com/r/Jokes/comments/4q0noj/why_does_superman_have_to_wait_until_tomorrow_to/,self.jokes,,He can't face the Crips tonight.,Why does Superman have to wait until tomorrow to fight gang violence in LA?,0
post,4q0ndb,2qh72,jokes,false,1466988369,https://old.reddit.com/r/Jokes/comments/4q0ndb/jaques_the_lumberjack_takes_a_barmaid_home_for/,self.jokes,,"Just outside a small town in Quebec lived a lumberjack by the name of Jacques. One day, as Jacques is done his work, he heads into the town as he normally does, and goes straight to the bar. He soon gets a few drinks in him, all the while, chatting up the barmaid. The barmaid is smitten by Jacques and agrees to go back to his place for the night.
After a passionate night with Jacques, the barmaid gets dressed the next morning, and heads out the door leaving Jacques to sleep in.
BANG! BANG! BANG!
Awoken by loud knocking on his door, Jacques jumps out of bed thinking the barmaid is back for more. To his surprise, two police officers stood at his door.
""What seems to be zee problem, officer?"" Jacques asks.
""It would seem that you have had sex without consent"" replies one of the officers.
""But zat is impossible!"" Jacques exclaims in disbelief.
""We're going to need you to come with us, as it is illegal to have sex without consent"" The other officer informs.
Jacques is awe struck, and says to the two officers, ""step in, look around, this whole place reeks of cunt scent!""",Jaques the Lumberjack takes a barmaid home for some fun...,0
post,4q0n9f,2qh72,jokes,false,1466988315,https://old.reddit.com/r/Jokes/comments/4q0n9f/how_do_you_make_a_goldfish_old/,self.jokes,,Take away the G.,How do you make a goldfish old?,15
post,4q0n7k,2qh72,jokes,false,1466988291,https://old.reddit.com/r/Jokes/comments/4q0n7k/my_exwife_is_like_a_tornado/,self.jokes,,"First she blows, then she sucks, then she took my house and dog.",My ex-wife is like a tornado,67
post,4q0mir,2qh72,jokes,false,1466988002,https://old.reddit.com/r/Jokes/comments/4q0mir/jenny_craig_shares_take_a_hit_following_brexit/,self.jokes,,Pounds are dropping fine without it,Jenny Craig shares take a hit following Brexit,0
post,4q0mc8,2qh72,jokes,false,1466987927,https://old.reddit.com/r/Jokes/comments/4q0mc8/what_if_netflix_had_a_dating_service/,self.jokes,,[deleted],What if Netflix had a dating service?,0
post,4q0m8s,2qh72,jokes,false,1466987885,https://old.reddit.com/r/Jokes/comments/4q0m8s/what_did_the_spring_peeper_frog_say_to_the_cow/,self.jokes,,Nice tits. ,What did the spring peeper (frog) say to the cow?,0
post,4q0m3n,2qh72,jokes,false,1466987818,https://old.reddit.com/r/Jokes/comments/4q0m3n/what_does_samuel_l_jackson_say_when_he_sees/,self.jokes,,[deleted],What does Samuel L. Jackson say when he sees people toss their used cigarettes on the street?,0
post,4q0jnq,2qh72,jokes,false,1466986833,https://old.reddit.com/r/Jokes/comments/4q0jnq/i_got_swole_by_eating_chinese_food/,self.jokes,,[deleted],I got swole by eating Chinese food,0
post,4q0jis,2qh72,jokes,false,1466986781,https://old.reddit.com/r/Jokes/comments/4q0jis/what_did_bill_say_to_hillary_after_sex/,self.jokes,,"""I'll be home in 20 minutes.""",What did Bill say to Hillary after sex?,1
post,4q0ilq,2qh72,jokes,false,1466986396,https://old.reddit.com/r/Jokes/comments/4q0ilq/why_is_their_always_lightning_in_france/,self.jokes,,"Obviously, since lightning takes the path of least resistance.",Why is their always lightning in France?,120
post,4q0gjo,2qh72,jokes,false,1466985566,https://old.reddit.com/r/Jokes/comments/4q0gjo/just_walked_by_a_senior_center_celebrating_pride/,self.jokes,,... It looked like they were having a gay old time,Just walked by a senior center celebrating pride...,5
post,4q0g1c,2qh72,jokes,false,1466985349,https://old.reddit.com/r/Jokes/comments/4q0g1c/red_pill_vs_blue_pill/,self.jokes,,"After reading just one post on each SubReddit, I realized that if I was an atheist I'd say a Male wrote the Old Testament, and a Female The New Testament... Or is it the other way around... Crap",Red Pill vs. Blue Pill,0
post,4q0fha,2qh72,jokes,false,1466985121,https://old.reddit.com/r/Jokes/comments/4q0fha/mexico_is_starting_to_build_a_wall/,self.jokes,,They're worried about the Americans crossing the border when Trump is elected. ,Mexico is starting to build a wall,9
post,4q0fgx,2qh72,jokes,false,1466985118,https://old.reddit.com/r/Jokes/comments/4q0fgx/why_did_the_lebanese_kid_go_to_school/,self.jokes,,[deleted],Why did the Lebanese kid go to school?,0
post,4q0ei3,2qh72,jokes,false,1466984738,https://old.reddit.com/r/Jokes/comments/4q0ei3/theres_a_woman_with_a_colostomy_bag/,self.jokes,,"Her boyfriend says he wants to fuck her in the pooper...

Which hole does he use?",There's a woman with a colostomy bag.,0
post,4q0e0x,2qh72,jokes,false,1466984539,https://old.reddit.com/r/Jokes/comments/4q0e0x/thatll_do_england_that_will_do_shrek/,self.jokes,,[removed],"""That'll do England that will do""- Shrek",1
post,4q0dps,2qh72,jokes,false,1466984417,https://old.reddit.com/r/Jokes/comments/4q0dps/whats_the_difference_between_luke_skywalker_and_a/,self.jokes,,Luke Skywalker eventually finds out who his father is.,What's the difference between Luke Skywalker and a black man?,32
post,4q0c9s,2qh72,jokes,false,1466983859,https://old.reddit.com/r/Jokes/comments/4q0c9s/people_from_the_uk_have_been_exercising_more/,self.jokes,,They've lost a few pounds.,People from the UK have been exercising more.,5
post,4q0c7d,2qh72,jokes,false,1466983834,https://old.reddit.com/r/Jokes/comments/4q0c7d/a_priestess_makes_me_make_a_promise/,self.jokes,,"She made me **swear** to never fucking swear.

",A priestess makes me make a promise,0
post,4q0c3w,2qh72,jokes,false,1466983793,https://old.reddit.com/r/Jokes/comments/4q0c3w/what_separates_man_from_animal/,self.jokes,,Divorce.,What separates man from animal?,7
post,4q0bq5,2qh72,jokes,false,1466983651,https://old.reddit.com/r/Jokes/comments/4q0bq5/oral_sex/,self.jokes,,"At this stage of our marriage, me and the wife only practice oral sex. Whenever we pass each other, we both say , 'fuck you.'",ORAL SEX,24
post,4q0bjb,2qh72,jokes,false,1466983583,https://old.reddit.com/r/Jokes/comments/4q0bjb/whats_the_difference_between_a_rundown_bus_stop/,self.jokes,,"One is just a crusty bus station, and the other is a busty crustacean!",What's the difference between a run-down bus stop and a big-breasted lobster?,3
post,4q0bfd,2qh72,jokes,false,1466983543,https://old.reddit.com/r/Jokes/comments/4q0bfd/what_do_you_get_when_you_cross_a_joke_with_a/,self.jokes,,[removed],What do you get when you cross a joke with a rhetorical question?,1
post,4q0ap8,2qh72,jokes,false,1466983244,https://old.reddit.com/r/Jokes/comments/4q0ap8/lawyers_get_robbed/,self.jokes,,[removed],Lawyers get robbed,1
post,4q0a00,2qh72,jokes,false,1466982952,https://old.reddit.com/r/Jokes/comments/4q0a00/what_is_the_most_popular_european_cuisine_in/,self.jokes,,Chichén Itzá,What is the most popular European cuisine in Mexico?,0
post,4q09z3,2qh72,jokes,false,1466982941,https://old.reddit.com/r/Jokes/comments/4q09z3/how_do_you_tell_the_difference_between_a_sunni/,self.jokes,,The Sunni's are the ones with the Shiite blown out of them.,How do you tell the difference between a Sunni and a Shiite Muslim?,0
post,4q09xy,2qh72,jokes,false,1466982927,https://old.reddit.com/r/Jokes/comments/4q09xy/what_kind_of_food_saps_a_man_will_to_live/,self.jokes,,Wedding cake,What kind of food saps a man will to live,0
post,4q0941,2qh72,jokes,false,1466982605,https://old.reddit.com/r/Jokes/comments/4q0941/a_grasshopper_walks_into_a_bar/,self.jokes,,"A grasshopper walks into a bar, and the bartender says, ""Hey, we have a drink named after you!""
The grasshopper looks surprised and asks, ""You have a drink named Steve?""",A grasshopper walks into a bar,16
post,4q0933,2qh72,jokes,false,1466982600,https://old.reddit.com/r/Jokes/comments/4q0933/british_women_and_british_cousine/,self.jokes,,[deleted],British women and british cousine,1
post,4q08x9,2qh72,jokes,false,1466982535,https://old.reddit.com/r/Jokes/comments/4q08x9/usain_bolt_sprints_into_a_metal_bar/,self.jokes,,[deleted],Usain Bolt sprints into a metal bar...,0
post,4q08t7,2qh72,jokes,false,1466982488,https://old.reddit.com/r/Jokes/comments/4q08t7/what_is_the_difference_between_snowmen_and/,self.jokes,,A: Snowballs.,What is the difference between snowmen and snowwomen?,2
post,4q089w,2qh72,jokes,false,1466982276,https://old.reddit.com/r/Jokes/comments/4q089w/how_do_you_starve_a_black_guy/,self.jokes,,[deleted],How do you starve a black guy?,0
post,4q07vd,2qh72,jokes,false,1466982126,https://old.reddit.com/r/Jokes/comments/4q07vd/a_black_man_walks_into_a_hotel/,self.jokes,,[removed],A black man walks into a hotel,0
post,4q07rr,2qh72,jokes,false,1466982087,https://old.reddit.com/r/Jokes/comments/4q07rr/got_into_an_accident_while_getting_road_head_the/,self.jokes,,[deleted],Got into an accident while getting road head the other day.,0
post,4q06qf,2qh72,jokes,false,1466981693,https://old.reddit.com/r/Jokes/comments/4q06qf/do_you_know_the_joke_about_a_group_of_people/,self.jokes,,It's just a punchline,Do you know the joke about a group of people waiting for fruit juice?,1
post,4q0658,2qh72,jokes,false,1466981472,https://old.reddit.com/r/Jokes/comments/4q0658/give_me_please/,self.jokes,,[removed],"Give me, please?",0
post,4q05h0,2qh72,jokes,false,1466981209,https://old.reddit.com/r/Jokes/comments/4q05h0/what_did_the_band_consisting_only_of_postmen_call/,self.jokes,,Vanmailen.,What did the band consisting only of postmen call itself?,0
post,4q05dw,2qh72,jokes,false,1466981173,https://old.reddit.com/r/Jokes/comments/4q05dw/david_cameron_i_cant_live/,self.jokes,,without EU,David Cameron: I can't live...,3
post,4q05bi,2qh72,jokes,false,1466981150,https://old.reddit.com/r/Jokes/comments/4q05bi/why_did_the_troll_cross_the_road/,self.jokes,,[removed],why did the troll cross the road,0
post,4q051h,2qh72,jokes,false,1466981041,https://old.reddit.com/r/Jokes/comments/4q051h/its_a_shame_what_happened_to_the_dolphinss_parents/,self.jokes,,I can't imagine being an Orfin ,It's a shame what happened to the Dolphins's parents......,6
post,4q04vz,2qh72,jokes,false,1466980979,https://old.reddit.com/r/Jokes/comments/4q04vz/crack_ya_ribs/,self.jokes,,[removed],Crack ya Ribs,1
post,4q04h1,2qh72,jokes,false,1466980827,https://old.reddit.com/r/Jokes/comments/4q04h1/will_was_killed_during_his_first_battle_with_the/,self.jokes,,"His comrades got confused when their commander yelled: ""Fire at Will!""",Will was killed during his first battle with the US army,4
post,4q04cx,2qh72,jokes,false,1466980781,https://old.reddit.com/r/Jokes/comments/4q04cx/an_englishman_a_scotsman_and_an_irishman_went_to/,self.jokes,,[deleted],"An Englishman, a Scotsman and an Irishman went to a bar.",1
post,4q03lp,2qh72,jokes,false,1466980495,https://old.reddit.com/r/Jokes/comments/4q03lp/knock_knock/,self.jokes,,"Who's there?

Alask.

Alask who? 

Alaska later",Knock Knock,1
post,4q02cp,2qh72,jokes,false,1466980008,https://old.reddit.com/r/Jokes/comments/4q02cp/what_do_you_call_the_reptile_that_started_the/,self.jokes,,The insti-gator. ,What do you call the reptile that started the fight?,7
post,4q022c,2qh72,jokes,false,1466979886,https://old.reddit.com/r/Jokes/comments/4q022c/a_coin_with_the_face_hillary_and_donald_on_each/,self.jokes,,[removed],"A coin with the face Hillary and Donald on each side. You flip it 319 million times, who loses??? Everyone!",2
post,4q01fs,2qh72,jokes,false,1466979636,https://old.reddit.com/r/Jokes/comments/4q01fs/i_like_my_love_like_i_like_my_cornbread/,self.jokes,,[deleted],I like my love like I like my cornbread...,0
post,4q018x,2qh72,jokes,false,1466979564,https://old.reddit.com/r/Jokes/comments/4q018x/why_did_the_cow_go_to_the_psychiatrist/,self.jokes,,[deleted],Why did the cow go to the psychiatrist?,0
post,4q00wf,2qh72,jokes,false,1466979422,https://old.reddit.com/r/Jokes/comments/4q00wf/a_tourist_goes_to_a_restaurant_in_spain/,self.jokes,,"and sees a pair of huge testicles on the counter. He asks the waiter what those are, and the waiter said, ""Today, there was a bullfight. These are the balls of the bull. You can eat them."" 

The man replied, ""I would like to!""

""Sorry,"" the waiter said, ""but these balls are already reserved for someone else. Come back tomorrow.""

The man does, and the waiter serves him his balls. However, they were very small! He gets angry at the waiter, and asks him about the testicles.

""Well, sometimes the bull wins.""",A tourist goes to a restaurant in Spain,27
post,4q00ig,2qh72,jokes,false,1466979282,https://old.reddit.com/r/Jokes/comments/4q00ig/how_much_space_does_the_eu_have_left/,self.jokes,,1GB,How much space does the EU have left?,0
post,4pzzop,2qh72,jokes,false,1466978957,https://old.reddit.com/r/Jokes/comments/4pzzop/a_man_from_cape_horn/,self.jokes,,"There once was a man from Cape Horn,

Who wished he had never been born.

And he wouldn't have been

if his father had seen

that the end of the rubber was torn.",A Man from Cape Horn,2
post,4pzz4q,2qh72,jokes,false,1466978731,https://old.reddit.com/r/Jokes/comments/4pzz4q/when_the_us_went_to_the_moon/,self.jokes,,"...they planted the American Flag. After all these years the radiation from the Sun will have bleached it completely white, so now if Aliens find it they are going to think the French were there first.",When the US went to the moon....,690
post,4pzye8,2qh72,jokes,false,1466978446,https://old.reddit.com/r/Jokes/comments/4pzye8/a_man_walks_into_a_zoo/,self.jokes,,[removed],A man walks into a zoo,1
post,4pzy6u,2qh72,jokes,false,1466978363,https://old.reddit.com/r/Jokes/comments/4pzy6u/harry_potter/,self.jokes,,"How did Harry get down from the hill?

Walking, jk rolling. ",Harry Potter,1
post,4pzxyx,2qh72,jokes,false,1466978272,https://old.reddit.com/r/Jokes/comments/4pzxyx/wanna_hear_a_racist_joke/,self.jokes,,Donald Trump.,Wanna hear a racist joke?,0
post,4pzxiy,2qh72,jokes,false,1466978106,https://old.reddit.com/r/Jokes/comments/4pzxiy/in_soviet_russia/,self.jokes,,...end of joke is when line punches *you*.,In Soviet Russia...,7
post,4pzw93,2qh72,jokes,false,1466977619,https://old.reddit.com/r/Jokes/comments/4pzw93/what_did_you_have_for_breakfast_pea_soup/,self.jokes,,"Q: What did you have for lunch?  
A: Pea Soup  
Q: What did you have for dinner?  
A: Pea Soup  
Q: What did you do all night?  
A: Pee soup…",What did you have for breakfast? Pea Soup,9
post,4pzw78,2qh72,jokes,false,1466977594,https://old.reddit.com/r/Jokes/comments/4pzw78/why_did_the_investment_bankers_start_dating/,self.jokes,,Compound interest,Why did the investment bankers start dating?,6
post,4pzw4d,2qh72,jokes,false,1466977564,https://old.reddit.com/r/Jokes/comments/4pzw4d/whats_invisible_and_smells_like_mice/,self.jokes,,Cat Farts...,What's Invisible and Smells Like Mice?,16
post,4pzvzd,2qh72,jokes,false,1466977503,https://old.reddit.com/r/Jokes/comments/4pzvzd/what_did_the_chemist_say_when_he_found_2_isotopes/,self.jokes,,HeHe ,What did the chemist say when he found 2 isotopes of helium?,38
post,4pzvw8,2qh72,jokes,false,1466977469,https://old.reddit.com/r/Jokes/comments/4pzvw8/what_do_you_get_a_german_child_for_his_birthday/,self.jokes,,[deleted],What do you get a German child for his birthday ?,0
post,4pzvsf,2qh72,jokes,false,1466977418,https://old.reddit.com/r/Jokes/comments/4pzvsf/what_do_you_call_a_25_year_old_male_who_plays/,self.jokes,,Single,What do you call a 25 year old male who plays Minecraft?,0
post,4pzvfj,2qh72,jokes,false,1466977282,https://old.reddit.com/r/Jokes/comments/4pzvfj/what_is_the_skinniest_animal/,self.jokes,,[deleted],What is the skinniest animal?,0
post,4pzv46,2qh72,jokes,false,1466977166,https://old.reddit.com/r/Jokes/comments/4pzv46/brexit_was_a_great_diet_plan/,self.jokes,,...because everyone in the UK lost a few pounds overnight.,Brexit was a great diet plan,1
post,4pzujb,2qh72,jokes,false,1466976963,https://old.reddit.com/r/Jokes/comments/4pzujb/an_eccentric_billionaire_throws_a_lavish_party/,self.jokes,,"Please bear with me as I heard/read this one years ago so I might not recall the details correctly:

An eccentric billionaire is throwing a lavish party with guests from all over the world. As the party is well under way he asks his guests to walk over to his Olympic sized swimming pool where he had it filled with all kinds of dangerous creatures, sharks, piranhas, crocodiles, you name it it is there! So he tells his guests ""I will give anything to the person who is brave enough to jump in the pool and swim across!"" The place falls silent as the guests only whisper amongst themselves in bewilderment. ""Anything that person can dream of will be his!"" the billionaire tells the guests again. Suddenly a large splash is heard and a guy is seen struggling to swim through, and miraculously he makes it across! The room erupts in cheers and the billionaire approaches the man who swam across, and tells him ""I am a man of my word, and since you made it across what do you desire? Money, mansions, my daughters hand in marriage?"" The man still visibly shaken and struggling to catch his breath replies ""I just want to know the name of the son of a bitch who pushed me in the pool!""
",An eccentric billionaire throws a lavish party...,65
post,4pzu6b,2qh72,jokes,false,1466976838,https://old.reddit.com/r/Jokes/comments/4pzu6b/an_american_pow_was_being_held_in_germany/,self.jokes,,"Both of his arms were injured during the fighting and the Nazis amputated one.

""Can you drop my arm over allied territory for my wife?"" The soldier asked. 

The doctors obliged. 
A few days later the other arm became infected and they amputated that one. 

""Can you drop it over allied territory for my wife?"" He asked again. 

The doctors met his second request. 

A few weeks later, the soldier's leg got smashed in the work camp and had to be amputated. 

""Can you drop my leg over allied territory for my wife?"" He asked. 

""Nein!"" The doctors told him. ""We cannot do this any more!""

""Why not?""

""We think you're  trying to escape!""






",An American POW was being held in Germany...,65
post,4pzu5d,2qh72,jokes,false,1466976831,https://old.reddit.com/r/Jokes/comments/4pzu5d/the_eu_is_much_like_a_bad_fart/,self.jokes,,Better out than in.,The EU is much like a bad fart.,2
post,4pztui,2qh72,jokes,false,1466976719,https://old.reddit.com/r/Jokes/comments/4pztui/a_girl_once_told_me_to_come_over_because_no_one/,self.jokes,,[deleted],A girl once told me to come over because no one was home,0
post,4pztcp,2qh72,jokes,false,1466976511,https://old.reddit.com/r/Jokes/comments/4pztcp/whats_the_difference_between_a_chick_pea_and_a/,self.jokes,,I've never had a lentil on my chest.,What's the difference between a chick pea and a lentil?,6
post,4pzt2d,2qh72,jokes,false,1466976405,https://old.reddit.com/r/Jokes/comments/4pzt2d/i_took_a_shit_today/,self.jokes,,[deleted],I took a shit today.,1
post,4pzsq0,2qh72,jokes,false,1466976268,https://old.reddit.com/r/Jokes/comments/4pzsq0/there_has_been_too_many_deaths_this_year/,self.jokes,,"
Like...

Alan Rickman

Anton Yelchin

Prince

Muhammad Ali

David Bowie

The UK",there has been too many deaths this year,0
post,4pzskz,2qh72,jokes,false,1466976215,https://old.reddit.com/r/Jokes/comments/4pzskz/nsfw_my_neighbors_favorite_body_organ_is_the/,self.jokes,,He's a pedophile with a patellar fetish.,[NSFW] My neighbor's favorite body organ is the kidney.,1
post,4pzsdy,2qh72,jokes,false,1466976139,https://old.reddit.com/r/Jokes/comments/4pzsdy/a_scottish_man_walks_store/,self.jokes,,"He asked for 15 litres of the best whiskey the clerk has. ""Did you bring a container for this?"" The clerk asks. ""You're speaking to it."" ",A Scottish man walks store...,12
post,4pzs4p,2qh72,jokes,false,1466976033,https://old.reddit.com/r/Jokes/comments/4pzs4p/what_do_you_call_a_joke_thats_about_people_dying/,self.jokes,,[deleted],What do you call a joke that's about people dying and nobody laughs at it?,0
post,4pzrze,2qh72,jokes,false,1466975978,https://old.reddit.com/r/Jokes/comments/4pzrze/the_eu_has_just_formed_a_new_dance_group/,self.jokes,,"It's called ""Free Movement"".",The EU has just formed a new dance group!,0
post,4pzr08,2qh72,jokes,false,1466975617,https://old.reddit.com/r/Jokes/comments/4pzr08/three_men_get_stranded_on_an_island/,self.jokes,,[deleted],Three men get stranded on an island.,0
post,4pzqxf,2qh72,jokes,false,1466975591,https://old.reddit.com/r/Jokes/comments/4pzqxf/an_american_a_brit_and_an_irishman_are_sitting_at/,self.jokes,,"A fly lands in each of their beers, the American takes the fly out of the glass and keeps on drinking. The Brit looks at the fly and asks the waitress for a new drink. The Irishman grabs the fly, squeezes it and yells ""spit it out you greedy bastard!""","An American, a Brit, and an Irishman are sitting at a bar",16
post,4pzqvm,2qh72,jokes,false,1466975573,https://old.reddit.com/r/Jokes/comments/4pzqvm/kelloggs_just_released_its_new_brexit_themed/,self.jokes,,[deleted],Kellogg's™ just released it's new Brexit themed waffles...,0
post,4pzpph,2qh72,jokes,false,1466975117,https://old.reddit.com/r/Jokes/comments/4pzpph/what_do_lebron_james_and_james_brown_have_in/,self.jokes,,They're both nicknamed the king and they both are overrated. ,What do Lebron James and James Brown have in common?,0
post,4pzpku,2qh72,jokes,false,1466975064,https://old.reddit.com/r/Jokes/comments/4pzpku/how_can_tell_if_theres_an_italian_at_the_cockfight/,self.jokes,,"He brings the duck

How can you tell if there's a Sicilian at the cockfight?

He bets on the duck

How can you tell if the Mafia is at the cockfight?

The duck wins",How can tell if there's an Italian at the cockfight?,4
post,4pzpiu,2qh72,jokes,false,1466975046,https://old.reddit.com/r/Jokes/comments/4pzpiu/a_philosopher_a_mathematician_and_an_idiot_were/,self.jokes,,"Suddenly, the three men found themselves standing before the pearly gates of Heaven, where St. Peter and the Devil were standing nearby.  

""Gentlemen,"" the Devil started, ""Due to the fact that Heaven is now overcrowded, St. Peter has agreed to limit the number of people entering Heaven. If anyone of you can ask me a question which I don't know or cannot answer, then you're worthy enough to go to Heaven; if not, then you'll come with me to Hell.""  

The philosopher then stepped up. 

""OK, give me the most comprehensive report on Socrates' teachings.""  

With a snap of his finger, a stack of paper appeared next to the Devil.  The philosopher read it and concluded it was correct. 

""Then go to hell!"" 

With another snap of his finger, the philosopher disappeared.  The mathematician then asked,

""Give me the most complicated formula ever theorized!"" 

With a snap of his finger, another stack of paper appeared next to the Devil. The mathematician read it and reluctantly agreed it was correct. 

""Then go to Hell!"" 

With another snap of his finger, the mathematician disappeared too.  The idiot then stepped forward and said, 

""Bring me a chair!""  

The Devil brought forward a chair. 

""Drill 7 holes on the seat."" 

The Devil did just that.  

The idiot then sat on the chair and let out a very loud fart.  Standing up, he asked, 

""Which hole did my fart come out from?""  

The Devil inspected the seat and said,

""The third hole from the right."" 

""Wrong,"" said the idiot, ""it's from my asshole.""  And the idiot went to heaven.","A philosopher, a mathematician and an idiot were riding in a car when it crashed into a tree.",119
post,4pzorr,2qh72,jokes,false,1466974770,https://old.reddit.com/r/Jokes/comments/4pzorr/britain_now_has_a_petition_to_void_the_eu/,self.jokes,,[deleted],"Britain now has a petition to void the EU referendum, and they called it...",2
post,4pzoa5,2qh72,jokes,false,1466974593,https://old.reddit.com/r/Jokes/comments/4pzoa5/some_people_think_its_difficult_to_live_with/,self.jokes,,"But really, it's not that hard.",Some people think it's difficult to live with Erectile Dysfunction,182
post,4pzna1,2qh72,jokes,false,1466974209,https://old.reddit.com/r/Jokes/comments/4pzna1/two_boys_were_arguing_when_the_teacher_entered/,self.jokes,,"Two boys were arguing when the teacher entered the room.

The teacher says, “Why are you arguing?”

One boy answers, “We found a ten dollor bill and decided to give it to whoever tells the biggest lie.”

“You should be ashamed of yourselves,” said the teacher, “When I was your age I didn’t even know what a lie was.”

The boys gave the ten dollars to the teacher.

IT HURTS!!!!!!!!!!!!!!!",Two boys were arguing when the teacher entered the room.,9
post,4pzn8e,2qh72,jokes,false,1466974191,https://old.reddit.com/r/Jokes/comments/4pzn8e/i_went_to_see_a_german_barber_and_said_can_i_have/,self.jokes,,"He said ""Yahs"", so I replied ""No, just the face.""","I went to see a German barber and said ""Can I have a shave please?""",0
post,4pzn21,2qh72,jokes,false,1466974130,https://old.reddit.com/r/Jokes/comments/4pzn21/a_guy_walks_into_a_bar/,self.jokes,,"He sees a pirate with a steering wheel in his pants. 

The guy asks ""Why do you have a steering wheel in your pants?"".

The pirate says ""I don't know but its driving me nuts!"".
",A guy walks into a bar.,5
post,4pzmjr,2qh72,jokes,false,1466973921,https://old.reddit.com/r/Jokes/comments/4pzmjr/a_man_with_no_job_no_family_no_money_and_every/,self.jokes,,"At the funeral, the eulogist said ""Wow his life sucked!""","A man with no job, no family, no money, and every cancer ever made got shot under the bridge he lived at because he was homeless",0
post,4pzkqo,2qh72,jokes,false,1466973244,https://old.reddit.com/r/Jokes/comments/4pzkqo/whats_worse_than_ten_children_in_one_bucket/,self.jokes,,One child in ten buckets.,What's worse than ten children in one bucket?,0
post,4pzk1t,2qh72,jokes,false,1466972997,https://old.reddit.com/r/Jokes/comments/4pzk1t/a_lumberjack_is_looking_for_work/,self.jokes,,[removed],A lumberjack is looking for work,1
post,4pzj5k,2qh72,jokes,false,1466972660,https://old.reddit.com/r/Jokes/comments/4pzj5k/what_do_you_call_a_group_of_black_researchers_on/,self.jokes,,A group of researchers you racist fuck. ,What do you call a group of black researchers on Antarctica?,0
post,4pzi8u,2qh72,jokes,false,1466972356,https://old.reddit.com/r/Jokes/comments/4pzi8u/i_opened_a_new_nightclub_named_erectile/,self.jokes,,"It was a complete flop, nobody came.",I opened a new nightclub named 'Erectile Dysfunction'.,11
post,4pzhum,2qh72,jokes,false,1466972205,https://old.reddit.com/r/Jokes/comments/4pzhum/a_man_goes_into_a_job_interview/,self.jokes,,"A man goes into a job interview, and presents himself well.

The employer is shocked at how professional he is, 

""Wow, you have an incredible resume, and present yourself fantastically, but you seem to be missing 5 years on this part of your resume. What happened there?""

The man replied ""Oh that's when I went to Yale.""

The employer is even more impressed. ""That's great, you're hired!""

The man is super happy and says ""Yay I got a yob!""",A man goes into a job interview...,574
post,4pzhsa,2qh72,jokes,false,1466972186,https://old.reddit.com/r/Jokes/comments/4pzhsa/a_guy_walks_into_a_store_to_try_to_find_a_suit/,self.jokes,,"A man is sitting in his house when he gets an invitation for his sister's wedding. However he doesn't own a suit.

So he heads down to the local suit store and asks the store owner if he has a suit for him.

""Yes I do!"" said the store owner, ""Right this way!""

The store owner leads the man through a row of purple suits, red suits, and green suits.

The man asks the store owner ""Don't you have any black suits?""

And the store owner replies to him ""No we didn't order any""",A guy walks into a store to try to find a suit for a wedding,0
post,4pzhlg,2qh72,jokes,false,1466972117,https://old.reddit.com/r/Jokes/comments/4pzhlg/yknow_i_hear_the_nword_a_hundred_times_a_day/,self.jokes,,I need to stop yelling it at black people.,Y'know I hear the N-word a hundred times a day...,4
post,4pzhex,2qh72,jokes,false,1466972055,https://old.reddit.com/r/Jokes/comments/4pzhex/why_dont_they_have_showers_on_airplanes/,self.jokes,,Because of the towel ban.,Why don't they have showers on airplanes?,26
post,4pzgd2,2qh72,jokes,false,1466971689,https://old.reddit.com/r/Jokes/comments/4pzgd2/two_guys_are_walking_their_dogs_down_the_street/,self.jokes,,"One has a golden retriever the other a Chihuahua. As they are going along the one with the retriever sees a bar. He turns to his friend and suggests they go in for a quick drink. His friend says ""That would be great but see the sign, no dogs allowed"". The guy turns to him and says ""Don't worry, just do what I do"". So the guy puts on some sunglasses and goes into the bar with his retriever. The tender turns to him and says ""Hey! No dogs allowed"". The guy quickly retorts ""Oh no, this is my seeing eye dog"". The bartender says ok and lets him sit.


His friend thinks about it and figures, why not. He puts on some sunglasses and walks in. The tender quickly turns and yells, ""Hey! No dogs allowed in the bar!""


The friend quickly replies ""No, you don't understand. This is my seeing eye dog!""


The bartender replies skeptically ""A Chihuahua is your seeing eye dog?""

""THEY GAVE ME A CHIHUAHUA?!""",Two guys are walking their dogs down the street...,285
post,4pzfet,2qh72,jokes,false,1466971354,https://old.reddit.com/r/Jokes/comments/4pzfet/a_professor_a_ceo_and_a_janitor_are_in_a_forest/,self.jokes,,"The fairy says ""I will give you what you most desire if you do someone else's job for a day.""

The professor says ""I'll be an elementary school teacher. What can be so hard about teaching a bunch of 6-year-olds how to read?"" so he is teleported into a classroom. After a few minutes, all the kids' screaming gets to his nerves, so he throws all his supplies and gives up.

The C.E.O says ""I'll be a waiter. All you do is carry food back and forth. This'll be a breeze"" so he is teleported to a restaurant. After about an hour, all the annoying customers drive him insane, so he smashes his plates on the ground and gives up.

The janitor says ""I'll be an artist"" so he is transported to an art facility. He glues all the classroom supplies and shattered plates to a canvas, then sells it for a billion dollars. The fairy asks the janitor how he was so clever.

The janitor says ""I got a masters degree in art.""","A professor, a CEO, and a janitor are in a forest when they discover a magic fairy.",1564
post,4pzfax,2qh72,jokes,false,1466971312,https://old.reddit.com/r/Jokes/comments/4pzfax/what_do_lawyers_call_hell/,self.jokes,,Home,What do lawyers call hell?,0
post,4pzevs,2qh72,jokes,false,1466971161,https://old.reddit.com/r/Jokes/comments/4pzevs/til_that_movie_bicycle_thieves_1948_didnt_had/,self.jokes,,That's racist!,"TIL that movie Bicycle Thieves (1948), didn't had black people in it...",0
post,4pzdr2,2qh72,jokes,false,1466970736,https://old.reddit.com/r/Jokes/comments/4pzdr2/how_do_you_stop_bacon_from_curling/,self.jokes,,You take away their brooms,How do you stop bacon from curling?,0
post,4pzdk9,2qh72,jokes,false,1466970665,https://old.reddit.com/r/Jokes/comments/4pzdk9/average_iq_of_the_eu_went_up/,self.jokes,,Thanks Brexit!,Average IQ of the EU went up,0
post,4pzdgc,2qh72,jokes,false,1466970628,https://old.reddit.com/r/Jokes/comments/4pzdgc/the_uk_summarized_in_two_sentences/,self.jokes,,"""No Scotland, you cannot leave the UK.""
""Hey Scotland, let's leave the EU.""",The U.K. Summarized in two sentences.,0
post,4pzbym,2qh72,jokes,false,1466970087,https://old.reddit.com/r/Jokes/comments/4pzbym/gay_bar_joke/,self.jokes,,[deleted],Gay bar joke,0
post,4pzb54,2qh72,jokes,false,1466969820,https://old.reddit.com/r/Jokes/comments/4pzb54/got_punched_in_the_face_by_a_convertible_car_the/,self.jokes,,...it's ruthless ,Got punched in the face by a convertible car the other day,0
post,4pzau6,2qh72,jokes,false,1466969719,https://old.reddit.com/r/Jokes/comments/4pzau6/a_novice_skier/,self.jokes,,Often jumps to contusions.,A Novice Skier,0
post,4pzagd,2qh72,jokes,false,1466969566,https://old.reddit.com/r/Jokes/comments/4pzagd/why_did_the_astronauts_abort_mission/,self.jokes,,[deleted],Why did the astronauts abort Mission?,0
post,4pza68,2qh72,jokes,false,1466969461,https://old.reddit.com/r/Jokes/comments/4pza68/all_day_ive_tried_to_convince_people_im_english/,self.jokes,,I'm leaving now,All day I've tried to convince people I'm English but I failed...,0
post,4pz9pr,2qh72,jokes,false,1466969310,https://old.reddit.com/r/Jokes/comments/4pz9pr/what_do_you_call_a_fish_with_no_eyes/,self.jokes,,Fsh,What do you call a fish with no eyes?,6
post,4pz9nm,2qh72,jokes,false,1466969289,https://old.reddit.com/r/Jokes/comments/4pz9nm/latvian_joke_q_what_are_one_potato_say_other/,self.jokes,,[removed],Latvian joke. •Q: What are one potato say other potato? •A: Premise stupid. Who have two potato?,1
post,4pz9bu,2qh72,jokes,false,1466969171,https://old.reddit.com/r/Jokes/comments/4pz9bu/what_do_you_call_a_field_used_to_grow_bows_and/,self.jokes,,An archerd.,What do you call a field used to grow bows and arrows?,0
post,4pz8pt,2qh72,jokes,false,1466968948,https://old.reddit.com/r/Jokes/comments/4pz8pt/why_is_santas_sack_so_big/,self.jokes,,[deleted],Why is Santa's sack so big?,12
post,4pz8nq,2qh72,jokes,false,1466968927,https://old.reddit.com/r/Jokes/comments/4pz8nq/i_was_playing_splat_zones_last_night/,self.jokes,,"An enemy squid was coming at me so I threw a Splash Wall to block him... But then I realized that I actually have Splat Bombs.

Edit: Whoops, wrong sub.",I was playing Splat Zones last night,0
post,4pz8f2,2qh72,jokes,false,1466968838,https://old.reddit.com/r/Jokes/comments/4pz8f2/you_really_have_to_hand_it_to_blind_prostitutes/,self.jokes,,[removed],You really have to hand it to blind prostitutes,1
post,4pz81o,2qh72,jokes,false,1466968700,https://old.reddit.com/r/Jokes/comments/4pz81o/how_was_the_copper_wire_invented/,self.jokes,,By two Jews who were fighting over a penny.,How was the copper wire invented?,0
post,4pz6wl,2qh72,jokes,false,1466968263,https://old.reddit.com/r/Jokes/comments/4pz6wl/the_owner_of_bell_incorporated_has_just_died/,self.jokes,,"The first in line to receive the inheritance is the owner's son, who gladly accepts it. However, the company lawyer says that he needs to take a photo of him for legal purposes. After developing the photo, he sends it off to the employees in the company to announce their new boss. He says ""Here's the fresh prints of Bell heir"".",The owner of Bell Incorporated has just died...,33
post,4pz6t1,2qh72,jokes,false,1466968234,https://old.reddit.com/r/Jokes/comments/4pz6t1/why_was_the_man_accused_of_sexual_harassment/,self.jokes,,He was a policeman,Why was the man accused of sexual harassment never arrested?,0
post,4pz5fv,2qh72,jokes,false,1466967753,https://old.reddit.com/r/Jokes/comments/4pz5fv/if_black_people_have_the_race_card_women_have_the/,self.jokes,,The Trump card.,"If black people have the race card, women have the gender card, what do rednecks have?",440
post,4pz4yz,2qh72,jokes,false,1466967587,https://old.reddit.com/r/Jokes/comments/4pz4yz/epicurean_oneliner/,self.jokes,,The epileptic eats burgers and shakes.,Epicurean One-Liner,0
post,4pz4rp,2qh72,jokes,false,1466967519,https://old.reddit.com/r/Jokes/comments/4pz4rp/the_captain_of_a_ship_got_into_a_fight_with_a_one/,self.jokes,,"Once the fight ended and he had prevailed he said to himself

""I lost a lot of good seamen today...""",The captain of a ship got into a fight with a one eyed monster...,0
post,4pz4ls,2qh72,jokes,false,1466967448,https://old.reddit.com/r/Jokes/comments/4pz4ls/a_pole_a_german_and_a_russian_go_to_prison/,self.jokes,,"A Pole, a German and a Russian are sent to prison. They each receive a 50-year sentence with no parole. The guard, when putting them in their cells, shows mercy on them and offers to give each of them a small supply of their favourite things to occupy their times. The Pole picks a collection of books by his favourite author, the German picks a case of strong beer, and the Russian picks a huge pack of cigarettes. After the 50 years pass, the guard checks on his prisoners. The Pole thanks the guard for allowing him to gain knowledge in his time, the German complains that he ran out of alcohol a week into his sentence, and the Russian asks the guard for a lighter.","A Pole, a German and a Russian go to prison...",271
post,4pz4cg,2qh72,jokes,false,1466967342,https://old.reddit.com/r/Jokes/comments/4pz4cg/how_can_you_tell_if_a_german_has_ocd/,self.jokes,,Ask them.  There's no other way.,How can you tell if a German has OCD?,0
post,4pz3er,2qh72,jokes,false,1466966988,https://old.reddit.com/r/Jokes/comments/4pz3er/in_the_middle_of_a_sermon_a_priest_openly/,self.jokes,,"After that, the congregation had a mass exodus.","In the middle of a sermon, a priest openly denounced the pope",0
post,4pz2q1,2qh72,jokes,false,1466966740,https://old.reddit.com/r/Jokes/comments/4pz2q1/whats_the_difference_between_a_cow_and_the/,self.jokes,,You can't milk a cow for 2000 years,What's the difference between a cow and the crucifixion?,6
post,4pz28e,2qh72,jokes,false,1466966545,https://old.reddit.com/r/Jokes/comments/4pz28e/what_do_you_call_an_indian_cowboy/,self.jokes,,Tex support,What do you call an Indian cowboy,1
post,4pz1g9,2qh72,jokes,false,1466966264,https://old.reddit.com/r/Jokes/comments/4pz1g9/my_mom_told_me_by_text_she_bought_me_a_box_of/,self.jokes,,[deleted],My mom told me by text she bought me a box of Gatorade,0
post,4pz0pw,2qh72,jokes,false,1466965989,https://old.reddit.com/r/Jokes/comments/4pz0pw/so_a_man_tries_to_buy_illegal_chicken_strips_at_a/,self.jokes,,[deleted],So a man tries to buy illegal chicken strips at a supermarket...,2
post,4pyzz8,2qh72,jokes,false,1466965713,https://old.reddit.com/r/Jokes/comments/4pyzz8/how_do_u_spell_candy_w_only_2_letters/,self.jokes,,c and y,How do u spell candy w only 2 letters,49
post,4pyziu,2qh72,jokes,false,1466965546,https://old.reddit.com/r/Jokes/comments/4pyziu/last_tuesday_i_farted/,self.jokes,,[removed],Last Tuesday I Farted.,0
post,4pyz50,2qh72,jokes,false,1466965401,https://old.reddit.com/r/Jokes/comments/4pyz50/2_niggers_walk_into_a_bar/,self.jokes,,[deleted],2 Niggers walk into a bar,0
post,4pyyqw,2qh72,jokes,false,1466965253,https://old.reddit.com/r/Jokes/comments/4pyyqw/i_love_the_new_snapchat_filters/,self.jokes,,[removed],I love the new snapchat filters...,1
post,4pyyed,2qh72,jokes,false,1466965119,https://old.reddit.com/r/Jokes/comments/4pyyed/what_is_jose_cuervos_favorite_book/,self.jokes,,Tequila Mockingbird.,What is Jose Cuervo's favorite book?,8
post,4pyybq,2qh72,jokes,false,1466965089,https://old.reddit.com/r/Jokes/comments/4pyybq/why_dont_bees_go_to_church/,self.jokes,,Because they are in sects.,Why don't bees go to church?,6
post,4pyxpx,2qh72,jokes,false,1466964846,https://old.reddit.com/r/Jokes/comments/4pyxpx/customer_feedback/,self.jokes,,"     A student at a management school came up to a pretty girl and hugged her without any warning.

The surprised girl said, “What was that?”

The guy smiled at her, “Direct marketing!”

The girl slapped him soundly.

“What was that?!” said the boy, holding his cheek.

      “Customer feedback.”
",“Customer feedback.”,22
post,4pyxf7,2qh72,jokes,false,1466964733,https://old.reddit.com/r/Jokes/comments/4pyxf7/there_are_a_lot_of_people_on_tinder_looking_for_a/,self.jokes,,"Honestly, tinder might be the absolute worst place to look for your missing friend. ","There are a lot of people on tinder ""looking for a friend""",0
post,4pyx21,2qh72,jokes,false,1466964577,https://old.reddit.com/r/Jokes/comments/4pyx21/president_obama_is_doing_his_morning_exercises/,self.jokes,,"...and jogging around the White House grounds when one of the Secret Service agents suggests he should see how fast he can circle the White House ten times. After all, it is a presidential tradition to try it at least once, and being moderately athletic, he figured he'd make pretty good time. So he stands at the south portico with the agent, who counts him down.

""3...2...1...go!""

President Obama takes off. He paces himself, not wanting to exhaust himself too quickly, and dodges gardeners, agents, and groundskeepers all the while. He laps the White House once, twice, three times, never losing speed. Several minutes pass by and as he laps the portico, the Secret Service agent yells out, ""One more, Mr. President!""

Obama launches himself into a mad sprint, going for broke and running like he'd never run before. He rounds one corner, then a second, then a third, and finally the last. Sweat is pouring down his face and his heart is pounding.

Finally, he reaches the portico and the agent clicks his stopwatch and hands Obama a cup of water. The president is very out of breath and bracing himself on the pillar, but pleased with himself all the same.

""So, how'd I do?""

The agent checks the stopwatch and says, ""Very well, Mr. President. Nine minutes and 23 seconds.""

""Really? That has to be a record!""

The agent responds, ""Not quite, sir. Bush did 9:11.""",President Obama is doing his morning exercises...,38
post,4pywkk,2qh72,jokes,false,1466964371,https://old.reddit.com/r/Jokes/comments/4pywkk/how_many_muslims_does_it_take_to_screw_in_a/,self.jokes,,Allah them,How many Muslims does it take to screw in a lightbulb?,32
post,4pyvzl,2qh72,jokes,false,1466964146,https://old.reddit.com/r/Jokes/comments/4pyvzl/a_man_walks_into_a_bar/,self.jokes,,[removed],A man walks into a bar.,0
post,4pyvz7,2qh72,jokes,false,1466964141,https://old.reddit.com/r/Jokes/comments/4pyvz7/fantastic_exercise/,self.jokes,,"Fantastic exercise that really helps you to lose weight: Turn your head to the left. Good. Turn your head to the right. Very good. Repeat this exercise whenever you are offered any food.

",Fantastic exercise,31
post,4pyvjp,2qh72,jokes,false,1466963975,https://old.reddit.com/r/Jokes/comments/4pyvjp/why_does_yoda_think_5_is_afraid_of_7/,self.jokes,,"Because ""6, 7 ate"".",Why does Yoda think 5 is afraid of 7?,1
post,4pyvja,2qh72,jokes,false,1466963969,https://old.reddit.com/r/Jokes/comments/4pyvja/whats_brown_smelly_and_sits_on_top_of_a_piano/,self.jokes,,Beethoven's last movement,"What's brown, smelly and sits on top of a piano?",1
post,4pyvco,2qh72,jokes,false,1466963896,https://old.reddit.com/r/Jokes/comments/4pyvco/once_my_mom_caught_me_conducting_lightning/,self.jokes,,...so she grounded me.,"Once, my mom caught me conducting lightning...",1
post,4pytz0,2qh72,jokes,false,1466963368,https://old.reddit.com/r/Jokes/comments/4pytz0/john_cena_payperview_matches_dont_sell_anymore_in/,self.jokes,,"Because when John Cena visits UK, EU can't see him.

*Ba dum tss*",John Cena pay-per-view matches don't sell anymore in the UK.,0
post,4pys50,2qh72,jokes,false,1466962678,https://old.reddit.com/r/Jokes/comments/4pys50/got_with_a_girl_for_the_first_time_last_night/,self.jokes,,[deleted],Got with a girl for the first time last night.,1
post,4pys0o,2qh72,jokes,false,1466962634,https://old.reddit.com/r/Jokes/comments/4pys0o/a_brand_new_cemetery_for_the_greats_now_will_let/,self.jokes,,Lots of people are dying to get in!,A brand new cemetery for the greats now will let anyone be buried there,0
post,4pyryq,2qh72,jokes,false,1466962608,https://old.reddit.com/r/Jokes/comments/4pyryq/teacher_did_your_father_help_your_with_your/,self.jokes,,[removed],Teacher: Did your father help your with your homework,1
post,4pyrws,2qh72,jokes,false,1466962587,https://old.reddit.com/r/Jokes/comments/4pyrws/an_old_man_on_his_deathbed_spent_his_entire_life/,self.jokes,,"Joke: An old man on his death bed has spent his entire life pinching pennies and clinging to all of his money. Friendless, he is surrounded by his priest, doctor, and lawyer. Just before he dies he tells them, ""I know most people say that you can't bring money with you after you die, but I want you to all throw this into my grave just as they are about to bury me."" With this being said he hands them all envelopes with $50,000 in them.

After his funeral the three are discussing the money. The doctor says, ""I have to confess something. I've really been wanting a vacation so I only threw $40,000 in.""

The priest follows, ""I must also confess. We are renovating the church so I only threw in $25,000. I feel terrible.""

The lawyer lashes out at them, ""You guys are terrible! Not only did I throw in the $50,000 he gave me, but I added my own $10,000.""

The doctor replies, ""Why in the world would you give that greedy man your money?""

The lawyer replies, ""He was a good man so I wrote him a check for the full amount.""",An old man on his deathbed spent his entire life clinging to his money,206
post,4pyrvv,2qh72,jokes,false,1466962577,https://old.reddit.com/r/Jokes/comments/4pyrvv/what_cereal_do_vote_leave_britains_eat/,self.jokes,,[removed],What cereal do vote leave Britains eat?,1
post,4pyrsk,2qh72,jokes,false,1466962546,https://old.reddit.com/r/Jokes/comments/4pyrsk/a_british_boy_and_his_grandfather_are_flying_to/,self.jokes,,"They pass over a city. The boy says ""Look, pap, aren't the city lights pretty?""

His grandfather answers ""I supposed, but I'm a tad disappointed.""

Confused, his grandson asks ""Why do you say that?""

His grandfather replies: ""Dresden isn't burning nearly as bright as it used to.""",A British boy and his grandfather are flying to Germany at night,1
post,4pyrad,2qh72,jokes,false,1466962340,https://old.reddit.com/r/Jokes/comments/4pyrad/a_polar_bears_wife_is_frustrated_with_her_bipolar/,self.jokes,,[deleted],A polar bear's wife is frustrated with her bipolar husband,0
post,4pyqdy,2qh72,jokes,false,1466962012,https://old.reddit.com/r/Jokes/comments/4pyqdy/how_do_you_recognize_a_limp_dick/,self.jokes,,He uses a crotch.,How do you recognize a limp dick?,0
post,4pyq5u,2qh72,jokes,false,1466961924,https://old.reddit.com/r/Jokes/comments/4pyq5u/gotta_admire_the_nazis_ethics_on_medical_research/,self.jokes,,...since they advanced the field without hurting any animals.,Gotta admire the Nazi's ethics on medical research...,2
post,4pyptm,2qh72,jokes,false,1466961785,https://old.reddit.com/r/Jokes/comments/4pyptm/i_call_my_friend_gator_because_he_likes_punching/,self.jokes,,He's a pecs predator.,I call my friend Gator because he likes punching people in the chest.,0
post,4pyprh,2qh72,jokes,false,1466961763,https://old.reddit.com/r/Jokes/comments/4pyprh/dirty_what_do_you_end_up_with_when_youre_too_lazy/,self.jokes,,[deleted],[Dirty] What do you end up with when you're too lazy to clean up after?,2
post,4pypo4,2qh72,jokes,false,1466961724,https://old.reddit.com/r/Jokes/comments/4pypo4/what_do_an_anorexic_girl_and_the_uk_have_in_common/,self.jokes,,They both lose pounds really fast.,What do an anorexic girl and the UK have in common?,41
post,4pyp4w,2qh72,jokes,false,1466961526,https://old.reddit.com/r/Jokes/comments/4pyp4w/whats_taylor_swifts_favorite_meal/,self.jokes,,[deleted],What's Taylor Swift's favorite meal?,0
post,4pyo35,2qh72,jokes,false,1466961100,https://old.reddit.com/r/Jokes/comments/4pyo35/when_australia_leaves_its_union/,self.jokes,,[deleted],When Australia leaves it's union....,0
post,4pymme,2qh72,jokes,false,1466960581,https://old.reddit.com/r/Jokes/comments/4pymme/so_i_went_to_visit_an_old_friend_with_a_stutter/,self.jokes,,"He had made quite a bit of money since we had seen each other and I asked him how he did it. ""Well I I go do door to do door and sel sell bibles"". I asked him how he had made so much doing it and he said that he just says ""yo you can b buy a bi bible or I I can re read iit to you"".",So I went to visit an old friend with a stutter...,12
post,4pymcs,2qh72,jokes,false,1466960484,https://old.reddit.com/r/Jokes/comments/4pymcs/what_was_the_problem_with_the_two_bears_who/,self.jokes,,[deleted],What was the problem with the two bears who played chess at the beach?,0
post,4pym8g,2qh72,jokes,false,1466960436,https://old.reddit.com/r/Jokes/comments/4pym8g/i_had_an_accident_today_at_the_ac_factory_i_work/,self.jokes,,[deleted],I had an accident today at the AC factory I work in.,8
post,4pym1j,2qh72,jokes,false,1466960368,https://old.reddit.com/r/Jokes/comments/4pym1j/trump_is_elected_president/,self.jokes,,And he finds out that he can't get anything done because of the USA's system of checks and balances.,Trump is elected president,0
post,4pylcz,2qh72,jokes,false,1466960092,https://old.reddit.com/r/Jokes/comments/4pylcz/my_old_classmate_became_a_nun/,self.jokes,,[deleted],My old classmate became a nun,0
post,4pykoy,2qh72,jokes,false,1466959821,https://old.reddit.com/r/Jokes/comments/4pykoy/not_safe_for_kids/,self.jokes,,Your parents are Santa clause AND the tooth fairy.,Not safe for kids,0
post,4pykl6,2qh72,jokes,false,1466959776,https://old.reddit.com/r/Jokes/comments/4pykl6/dirty_my_friend_has_a_pc/,self.jokes,,[deleted],[dirty] my friend has a pc,0
post,4pykfb,2qh72,jokes,false,1466959719,https://old.reddit.com/r/Jokes/comments/4pykfb/while_playing_in_the_backyard_johnny_kills_a/,self.jokes,,"While playing in the backyard, Little Johnny kills a honeybee. His father sees him killing the honeybee and angrily says, ""No honey for you for one month!"" Later that afternoon, Johnny's dad catches him tearing the wings off a butterfly. ""That's it! No butter for you for one month!"" says his dad. Later that evening as Johnny's mother cooks dinner, a cockroach run across the kitchen floor. She jumps and stomps on it, and then looks up to find Little Johnny and her husband watching her. Little Johnny looks at his father and says, ""Are you going to tell her, Dad, or do you want me to?","While playing in the backyard, Johnny kills a honeybee",77
post,4pyk79,2qh72,jokes,false,1466959623,https://old.reddit.com/r/Jokes/comments/4pyk79/a_village_kid_asks_his_parish_priest_if_he_could/,self.jokes,,"Priest: ""Ok but my horse is no ordinary horse. You have to pay attention to the instructions:
Say THANK GOD and it will bolt &amp; run. Say PRAISE YOU LORD &amp; it will run faster. Say LORD HAVE MERCY and it will stop immediately. Don't forget.""

So, the kid gets on the horse, says ""THANK GOD"" and they run off. Wanting to see how fast the horse can run, he says ""PRAISE YOU LORD"" repeatedly and the horse ran so fast, the kid didn't see that they were headed for a cliff. Alarmed, he wanted to stop but he couldn't remember the command. Just when they were about to fall off, he remembered &amp; exclaimed ""LORD HAVE MERCY!!!"". Instantly, the horse stopped just a few inches away from the edge.

Kid:"" Oh my god...jeez. boy, that was sooo close. whew! thank god!""",A village kid asks his parish priest if he could play with his horse..,16
post,4pyjey,2qh72,jokes,false,1466959285,https://old.reddit.com/r/Jokes/comments/4pyjey/what_do_you_call_4_mexicans_in_quicksand/,self.jokes,,"quatro cinco
",What do you call 4 Mexicans in quicksand?,11
post,4pyjb4,2qh72,jokes,false,1466959244,https://old.reddit.com/r/Jokes/comments/4pyjb4/whats_the_difference_between_a_pilsner_and_a_lager/,self.jokes,,I don't know any hipsters that try to dress like pilsners.,what's the difference between a pilsner and a lager?,0
post,4pyjat,2qh72,jokes,false,1466959241,https://old.reddit.com/r/Jokes/comments/4pyjat/a_drunk_walks_out_of_a_bar_one_morning/,self.jokes,,"He bumps into a cop.  The cop points at the bar and says, ""Hey, your eyes are all bloodshot, have you been drinking Bloody Marys in there?""  The drunk points to his cop car and says, ""Hey, your eyes are all glazed over, have you been eating donuts in there?""",A drunk walks out of a bar one morning...,2
post,4pyiyf,2qh72,jokes,false,1466959103,https://old.reddit.com/r/Jokes/comments/4pyiyf/a_little_boy_gets_on_the_public_bus_and_sits/,self.jokes,,"A little boy gets on the public bus and sits right behind the bus driver. The boy keeps repeatedly saying,"" If my mom was a cow and my dad was a bull, I'd be a little calf. If my mom was a hen and my dad was a chicken, I'd be a little chick. If my mom was a deer and my dad was a buck, I'd be a little deer. If my mom was a duck and my dad was a goose, I'd be a little duckling."" The bus annoyed bus driver stops the bus and turns to the boy saying, ""What if your mom was a drunk and you dad was a bum?"" The boy responds, ""Then I'd be a bus driver.""",A little boy gets on the public bus and sits right behind the bus driver,59
post,4pyis9,2qh72,jokes,false,1466959048,https://old.reddit.com/r/Jokes/comments/4pyis9/powerful_lost_love_spell_voodoo_spell_traditional/,self.jokes,,[removed],Powerful Lost Love spell Voodoo spell Traditional Healer +27633809460 @,1
post,4pyi6f,2qh72,jokes,false,1466958820,https://old.reddit.com/r/Jokes/comments/4pyi6f/job_application/,self.jokes,,"Apparently this is an actual job application submitted by a 17 year old boy at a McDonald's establishment in Florida... 

NAME: Greg Bulmash 

SEX: Not yet. Still waiting for the right person. 

DESIRED POSITION: Company's President or Vice President. But seriously, whatever's available. If I was in a position to be picky, I wouldn't be applying here in the first place. 

DESIRED SALARY: $185,000 a year plus stock options and a Michael Ovitz style severance package. If that's not possible, make an offer and we can haggle. 

EDUCATION: Yes. 

LAST POSITION HELD: Target for middle management hostility. 

SALARY: Less than I'm worth. 

MOST NOTABLE ACHIEVEMENT: My incredible collection of stolen pens and post-it notes. 

REASON FOR LEAVING: It sucked. 

HOURS AVAILABLE TO WORK: Any. 

PREFERRED HOURS: 1:30-3:30 p.m., Monday, Tuesday, and Thursday. 

DO YOU HAVE ANY SPECIAL SKILLS?: Yes, but they're better suited to a more intimate environment. 

MAY WE CONTACT YOUR CURRENT EMPLOYER?: If I had one, would I be here? 

DO YOU HAVE ANY PHYSICAL CONDITIONS THAT WOULD PROHIBIT YOU FROM LIFTING UP TO 50 LBS?: Of what? 

DO YOU HAVE A CAR?: I think the more appropriate question here would be ""Do you have a car that runs?"" 

HAVE YOU RECEIVED ANY SPECIAL AWARDS OR RECOGNITION?: I may already be a winner of the Publishers Clearing house Sweepstakes. 

DO YOU SMOKE?: On the job no, on my breaks yes. 

WHAT WOULD YOU LIKE TO BE DOING IN FIVE YEARS?: Living in the Bahamas with a fabulously wealthy dumb sexy blonde super model who thinks I'm the greatest thing since sliced bread. Actually, I'd like to be doing that now. 

DO YOU CERTIFY THAT THE ABOVE IS TRUE AND COMPLETE TO THE BEST OF YOUR KNOWLEDGE?: Yes. Absolutely. 

SIGN HERE: Aries.
",Job Application,119
post,4pyg7h,2qh72,jokes,false,1466958116,https://old.reddit.com/r/Jokes/comments/4pyg7h/why_do_people_who_drink_milk_struggle_to_walk/,self.jokes,,Because they lactose.,Why do people who drink milk struggle to walk?,28
post,4pydne,2qh72,jokes,false,1466957122,https://old.reddit.com/r/Jokes/comments/4pydne/how_long_does_it_take_a_group_of_mexicans_to/,self.jokes,,"Oh look, they're done. ",How long does it take a group of Mexicans to build a building?,1
post,4pyd9l,2qh72,jokes,false,1466956972,https://old.reddit.com/r/Jokes/comments/4pyd9l/what_do_you_call_a_faucet_that_wont_give_water_to/,self.jokes,,A sbigot.,What do you call a faucet that won't give water to gay people?,17
post,4pyc5w,2qh72,jokes,false,1466956536,https://old.reddit.com/r/Jokes/comments/4pyc5w/whats_the_deal_with_airline_peanuts/,self.jokes,,[removed],What's the deal with airline peanuts?,1
post,4pyb0k,2qh72,jokes,false,1466956087,https://old.reddit.com/r/Jokes/comments/4pyb0k/the_evening_news/,self.jokes,,"The evening news is the only place where they say ""Good Evening""  then proceed to tell you why it isn't.",The Evening News,18
post,4pyawr,2qh72,jokes,false,1466956047,https://old.reddit.com/r/Jokes/comments/4pyawr/why_did_everyone_disregard_the_midgets_stand_up/,self.jokes,,Because puns are the lowest form of comedy.,Why did everyone disregard the midget's stand up routine?,2
post,4pya3a,2qh72,jokes,false,1466955737,https://old.reddit.com/r/Jokes/comments/4pya3a/fuck_cheesy_chatup_lines_we_need_better_breakup/,self.jokes,,[deleted],"Fuck cheesy chat-up lines, we need better break-up lines:",0
post,4py9wi,2qh72,jokes,false,1466955663,https://old.reddit.com/r/Jokes/comments/4py9wi/a_depressed_monkey_wanted_to_end_his_life/,self.jokes,,[deleted],A depressed monkey wanted to end his life.,0
post,4py9ue,2qh72,jokes,false,1466955640,https://old.reddit.com/r/Jokes/comments/4py9ue/the_average_eu_woman_just_got_hotter/,self.jokes,,[removed],The average EU woman just got hotter,9653
post,4py9dc,2qh72,jokes,false,1466955447,https://old.reddit.com/r/Jokes/comments/4py9dc/there_is_no_such_thing_as_a_bad_joke/,self.jokes,,Only jokes with Jews and without.,There is no such thing as a bad joke,0
post,4py8fp,2qh72,jokes,false,1466955081,https://old.reddit.com/r/Jokes/comments/4py8fp/whats_a_mostly_red_rainbow_called/,self.jokes,,A pride flag found at Orlando.,What's a mostly red rainbow called?,0
post,4py86u,2qh72,jokes,false,1466954989,https://old.reddit.com/r/Jokes/comments/4py86u/whats_the_difference_between_a_seagull_and_a_baby/,self.jokes,,[deleted],What's the difference between a seagull and a baby?,1
post,4py86c,2qh72,jokes,false,1466954982,https://old.reddit.com/r/Jokes/comments/4py86c/how_many_police_officers_does_it_take_to_screw_in/,self.jokes,,"None, they just beat the shit out of the room for being black. ",How many police officers does it take to screw in a lightbulb?,0
post,4py83q,2qh72,jokes,false,1466954951,https://old.reddit.com/r/Jokes/comments/4py83q/a_man_is_stopped_for_speeding_on_the_highway/,self.jokes,,"The driver, when confronted by the cop to be issued a ticket, suddenly confesses that he has heroin with him in the vehicle.
Shocked, the cop calls for backup, explaining that the man who he caught speeding admitted that he had drugs on him.

A narcotics team arrives and searches the vehicle to find nothing of interest. Confronting the driver, they ask for an explanation. 

""The cop said I had heroin in my car?! Of course not!"" exclaims the driver. 

""I bet he told you I was speeding too""
",A man is stopped for speeding on the highway,110
post,4py83n,2qh72,jokes,false,1466954951,https://old.reddit.com/r/Jokes/comments/4py83n/news_headline_2016_glorious_victory_for_the_leave/,self.jokes,,"News headline 2116: UNITED EARTH SPACESHIP CRASHES ON THE BIG ISLAND OFF THE COAST OF EURASIA. ANGRY LOCAL TRIBESPEOPLE SACRIFICE CREW, EAT BRAINS",News headline 2016: GLORIOUS VICTORY FOR THE LEAVE CAMPAIGN. BRITAIN TO LEAVE THE EU,0
post,4py7vb,2qh72,jokes,false,1466954859,https://old.reddit.com/r/Jokes/comments/4py7vb/ad_for_a_wife/,self.jokes,,"A man inserted an 'ad' in the classifieds: ""Wife wanted.""  Next day he received a hundred letters.  They all said the same thing: ""You can have mine.""",ad for a wife,16
post,4py6z4,2qh72,jokes,false,1466954520,https://old.reddit.com/r/Jokes/comments/4py6z4/what_do_you_call_a_prostitute_with_a_runny_nose/,self.jokes,,Full,What do you call a prostitute with a runny nose?,60
post,4py6k1,2qh72,jokes,false,1466954360,https://old.reddit.com/r/Jokes/comments/4py6k1/why_did_dwayne_the_rock_johnson_have_to_change/,self.jokes,,"Because his nutritionist said he had too many minerals in his system!
","Why did Dwayne ""The Rock"" Johnson have to change his diet?",2
post,4py62o,2qh72,jokes,false,1466954158,https://old.reddit.com/r/Jokes/comments/4py62o/800_owed/,self.jokes,,"A man is getting into the shower just as his wife is finishing up her shower, when the doorbell rings. The wife quickly wraps herself in a towel and runs downstairs.  When she opens the door, there stands Bob, the next-door neighbor.  Before she says a word, Bob says, ""I’ll give you $800 to drop that towel.""  After thinking for a moment, the woman drops her towel and stands naked in front of Bob.  After a few seconds, Bob hands her $800 and leaves.  The woman wraps back up in the towel and goes back upstairs.  When she gets to the bathroom, her husband asks, ""Who was that?"" ""It was Bob the next door neighbor,"" she replies.  ""Great,"" the husband says, ""did he say anything about the $800 he owes me?"" ",$800 owed,57
post,4py5ws,2qh72,jokes,false,1466954107,https://old.reddit.com/r/Jokes/comments/4py5ws/when_kim_kardashian_is_off_camera_she_is_helping/,self.jokes,,Too bad she is always on camera. ,When Kim Kardashian is off camera she is helping little homeless kids.,1
post,4py5wk,2qh72,jokes,false,1466954106,https://old.reddit.com/r/Jokes/comments/4py5wk/emmanuel_lubezki_walks_into_a_bar/,self.jokes,,and orders one shot.,Emmanuel Lubezki walks into a bar,1
post,4py5u5,2qh72,jokes,false,1466954086,https://old.reddit.com/r/Jokes/comments/4py5u5/why_does_britain_like_tea_so_much/,self.jokes,,Because tea leaves.,Why does Britain like tea so much?,5540
post,4py5ib,2qh72,jokes,false,1466953967,https://old.reddit.com/r/Jokes/comments/4py5ib/marriage_the_real_story/,self.jokes,,"A husband walks into the bedroom to see his wife packing a suitcase. He asks, ""What are you doing?""
She answers, ""I'm moving to Nevada . I heard that prostitutes there get paid $400.00 for what I'm doing for YOU for FREE!""
Later that night, on her way out, the wife walks into the bedroom and sees her husband packing his suitcase.
When she asks him where he's going, he replies,
""I'm coming too. I want to see how you live on $800.00 a year.""","Marriage, the real story",364
post,4py5i4,2qh72,jokes,false,1466953965,https://old.reddit.com/r/Jokes/comments/4py5i4/how_do_you_start_a_stampede/,self.jokes,,"Go to a reddit meetup and yell ""Feminist!""",How do you start a stampede?,4
post,4py5c8,2qh72,jokes,false,1466953906,https://old.reddit.com/r/Jokes/comments/4py5c8/an_engineer_dies_and_goes_to_heaven/,self.jokes,,"He meets St. Peter at the pearly gates, and St. Peter checks the list. St. Peter doesn't find his name, so he says 'sorry, looks like you are supposed to go to the other place'.

So the engineer then goes down to Hell. Soon, he starts seeing things that could be improved. He builds a central air conditioning unit to help control the heat. He starts installing a central sewage system.

God notices, and quickly calls Satan. He calls and says 'there's been a mistake! The engineer is supposed to be up here with us!'

Satan replies: 'you know, we're pretty happy with what the changes he had been making, I think we'll keep him'

God gets mad and says 'you send him up here this minute or else I'll sue you!'

Satan laughs and says, 'yeah, you and what lawyers?'",An engineer dies and goes to heaven...,1231
post,4py56m,2qh72,jokes,false,1466953850,https://old.reddit.com/r/Jokes/comments/4py56m/pedophiles_are_fucking_immature_assholes/,self.jokes,,[removed],Pedophiles are fucking immature assholes,2
post,4py50s,2qh72,jokes,false,1466953790,https://old.reddit.com/r/Jokes/comments/4py50s/what_do_you_call_a_black_guy_in_outer_space/,self.jokes,,An astronaut you racist bastard. ,What do you call a black guy in outer space?,114
post,4py4zx,2qh72,jokes,false,1466953781,https://old.reddit.com/r/Jokes/comments/4py4zx/whats_the_difference_between_a_garbanzo_bean_and/,self.jokes,,I've never paid 200 dollars to have a garbanzo bean on my chest. ,What's the difference between a garbanzo bean and a chickpea?,6
post,4py4cd,2qh72,jokes,false,1466953542,https://old.reddit.com/r/Jokes/comments/4py4cd/while_its_technically_correct_that_muslims_have/,self.jokes,, they still only get one girl apiece. ,While it's technically correct that muslims have 72 virgins waiting for them in heaven...,0
post,4py414,2qh72,jokes,false,1466953415,https://old.reddit.com/r/Jokes/comments/4py414/there_is_a_chair/,self.jokes,,[deleted],There is a chair,0
post,4py3rh,2qh72,jokes,false,1466953302,https://old.reddit.com/r/Jokes/comments/4py3rh/whats_the_difference_between_a_lawyer_and_a/,self.jokes,,"One you pay $500 an hour to screw you.

The other one has sex for money.",What's the difference between a lawyer and a prostitute?,31
post,4py3pz,2qh72,jokes,false,1466953286,https://old.reddit.com/r/Jokes/comments/4py3pz/my_girlfriend_complained_about_my_obsession_with/,self.jokes,,"So I said, ""Bae, leave.""",My girlfriend complained about my obsession with spices.,19
post,4py30h,2qh72,jokes,false,1466952993,https://old.reddit.com/r/Jokes/comments/4py30h/whats_the_difference_between_a_garbanzo_beans_and/,self.jokes,,[deleted],What's the difference between a garbanzo beans and chickpea?,1
post,4py18l,2qh72,jokes,false,1466952239,https://old.reddit.com/r/Jokes/comments/4py18l/so_i_have_a_joke_about_pizza/,self.jokes,,...but it's too cheesy,So I have a joke about pizza...,15
post,4py16w,2qh72,jokes,false,1466952219,https://old.reddit.com/r/Jokes/comments/4py16w/now_that_britain_has_left_the_eu_youll_need_a/,self.jokes,,"...for everything else, there's Mastercard.","Now that Britain has left the EU, you'll need a Visa to get in and around",2
post,4py0sh,2qh72,jokes,false,1466952060,https://old.reddit.com/r/Jokes/comments/4py0sh/a_native_american_emerges_with_a_new_born/,self.jokes,,"A Native American chief emerges from a teepee with a new born in his hands, looks round at the crowd of awaiting people and announces, ""this boy shall be known as ""Sitting Bull"""". 

One young man approaches the chief and asks ""Chief, why name the boy ""Sitting Bull?""  

""It is simple. When I emerge from the teepee with a new born, I name him after the first thing I see. Like when I named your father. I emerged from teepee and saw the majestic sun rise, and so I named him ""Rising Sun"". Then with your brother, I emerge and see the moon glowing in the sky, so I name him ""Glowing Moon"". And just now, I emerge and see bull resting in field, so I name him ""Sitting Bull"". 

Why do you ask, Two Dogs Fucking?""",A Native American emerges with a new born...,11
post,4py0ln,2qh72,jokes,false,1466951984,https://old.reddit.com/r/Jokes/comments/4py0ln/hillary_clinton_doesnt_negotiate_with_countries/,self.jokes,,[deleted],Hillary Clinton doesn't negotiate with countries that sponsor terrorism...,15
post,4pxzvl,2qh72,jokes,false,1466951707,https://old.reddit.com/r/Jokes/comments/4pxzvl/what_did_the_japanese_man_say_as_the_hiroshima/,self.jokes,,Wow this blew up fast.,"What did the Japanese man say as the Hiroshima sky was filled with the light of an atomic bomb, in a split second?",10
post,4pxyqf,2qh72,jokes,false,1466951247,https://old.reddit.com/r/Jokes/comments/4pxyqf/what_did_the_metal_say_to_the_hydraulic_press/,self.jokes,,"""I'm impressed""",What did the metal say to the hydraulic press?,3
post,4pxwn7,2qh72,jokes,false,1466950329,https://old.reddit.com/r/Jokes/comments/4pxwn7/there_were_three_pows_together_in_a_british/,self.jokes,,"The British began by torturing the German. After long hours of silence infected by bloodcurdling screams, he talked, and was sent back to the prison, ashamed. He told the others what he had done and urged them to be stronger than he was.

They next began torturing the Japanese man. Through all the pain and agony, he stayed strong for three days, but in the end, talked. He was sent back to the prison, having brought shame to himself, his family, and his country.

They finally sent in the Italian. For an unending three weeks, they tortured him, until they realized if they did anything else to the poor man, he would die, so they sent him back. When he got back to the prison cell bloody and battered, the other POWs asked him, ""So? Did you talk?""

""How could I talk with my hands tied behind my back?""","There were three POWs together in a British prison in the Second World War, a German, a Japanese, and an Italian.",17966
post,4pxwl9,2qh72,jokes,false,1466950302,https://old.reddit.com/r/Jokes/comments/4pxwl9/a_man_walks_by_an_insane_asylum/,self.jokes,,"An man walks by an insane asylum and hears the inmates gleefully shouting ""21! 21! 21"" As he gets closer he sees a hole in the brick wall which he approaches so he can peek in and see what's going on. The inmates poke a stick through the hole, poking him in the eye, and yell ""22! 22! 22!""",A man walks by an insane asylum...,41
post,4pxwci,2qh72,jokes,false,1466950190,https://old.reddit.com/r/Jokes/comments/4pxwci/ive_spent_all_day_trying_to_convince_people_on/,self.jokes,,I give up.,I've spent all day trying to convince people on Reddit I'm French.,701
post,4pxvk3,2qh72,jokes,false,1466949842,https://old.reddit.com/r/Jokes/comments/4pxvk3/the_reason_i_dont_go_swimming_in_public_swimming/,self.jokes,,[removed],The reason I dont go swimming in public swimming pools is because of the alarming pH levels. It's almost all pee no H,1
post,4pxvc6,2qh72,jokes,false,1466949746,https://old.reddit.com/r/Jokes/comments/4pxvc6/some_kind_redditor_gave_me_gold/,self.jokes,,"it was AUmazing!

EDIT: AUsome! Someone just actually gilded this! THANK YOU!

EDIT2: AU no. He/She/It just took it back.",Some kind redditor gave me gold...,0
post,4pxt8q,2qh72,jokes,false,1466948787,https://old.reddit.com/r/Jokes/comments/4pxt8q/hyderabadi_whatsapp_joke/,self.jokes,,[removed],Hyderabadi whatsapp joke,1
post,4pxrhp,2qh72,jokes,false,1466947947,https://old.reddit.com/r/Jokes/comments/4pxrhp/did_you_hear_about_the_dyslexic_agnostic_insomniac/,self.jokes,,He stayed awake all night wondering if there really is a dog.,"Did you hear about the dyslexic, agnostic insomniac?",44
post,4pxrdz,2qh72,jokes,false,1466947903,https://old.reddit.com/r/Jokes/comments/4pxrdz/three_friends_decided_to_go_hunting_together/,self.jokes,,"One was a lawyer, one a doctor, and the other a preacher. As they were walking, along came a big buck. The three of them shot at the same time and the buck dropped immediately. The hunting party rushed to see how big it actually was. Upon reaching the fallen deer, they found out that it was dead but only had one bullet hole. A debate followed concerning whose buck it was. When a game warden came by, he offered to help. A few moments later, he had the answer. He said with much confidence, ""The pastor shot the buck!"" The friends were amazed that he could determine that so quickly and with so little examination. The game warden just smiled. ""It was easy to figure out. The bullet went in one ear and out the other.""",Three friends decided to go hunting together.,24
post,4pxr46,2qh72,jokes,false,1466947766,https://old.reddit.com/r/Jokes/comments/4pxr46/in_tesco_earlier_the_cashier_asked_the_foreign/,self.jokes,,"Fook me, we only voted out 2 days ago, give them a chance!!!","In Tesco earlier, the cashier asked the Foreign couple in front of me if they wanted help packing their bags.",2
post,4pxqxz,2qh72,jokes,false,1466947681,https://old.reddit.com/r/Jokes/comments/4pxqxz/a_blind_man_walks_past_the_fish_market_in_the/,self.jokes,,"and he says ""Good morning ladies"".",A blind man walks past the fish market in the morning,0
post,4pxqwe,2qh72,jokes,false,1466947663,https://old.reddit.com/r/Jokes/comments/4pxqwe/why_old_men_dont_get_hired/,self.jokes,,"An old man is before a human resource manager for a job interview.
The interviewer asks, ""What is your greatest weakness?"" The old man replies, ""Honesty."" The interviewer says, ""I don't think honesty is a weakness.""  The old man replies, ""I don't give a fuck what you think!""",Why old men don't get hired.,1
post,4pxqom,2qh72,jokes,false,1466947554,https://old.reddit.com/r/Jokes/comments/4pxqom/donald_trump_becomes_the_new_president/,self.jokes,,Yeah that's it. ,Donald Trump becomes the new president.,0
post,4pxq8e,2qh72,jokes,false,1466947318,https://old.reddit.com/r/Jokes/comments/4pxq8e/whats_the_worst_part_about_doing_crossfit/,self.jokes,,Having to shop at Kid's GAP. ,What's the worst part about doing crossfit?,5
post,4pxppf,2qh72,jokes,false,1466947075,https://old.reddit.com/r/Jokes/comments/4pxppf/how_many_gears_does_a_french_army_tank_have/,self.jokes,,[deleted],How many gears does a french army tank have?,1
post,4pxpja,2qh72,jokes,false,1466946990,https://old.reddit.com/r/Jokes/comments/4pxpja/what_disease_did_ben_and_jerry_give_to_all_of_the/,self.jokes,,[deleted],What disease did Ben and Jerry give to all of the prostitutes in Vermont?,0
post,4pxmel,2qh72,jokes,false,1466945387,https://old.reddit.com/r/Jokes/comments/4pxmel/a_trump_supporter_a_mexican_and_an_asian_person/,self.jokes,,"The pilot says that they need to throw out something that they already have a lot of.
The Mexican throws out a bag of tortillas, the Asian person throws out a bag of rice, and the Trump supporter throws out the Mexican.","A trump supporter, a Mexican, and an Asian person are on a plane when it starts going down",0
post,4pxmd0,2qh72,jokes,false,1466945363,https://old.reddit.com/r/Jokes/comments/4pxmd0/did_you_see_the_sun_had_an_exclusive_interview/,self.jokes,,[deleted],Did you see The Sun had an exclusive interview with Dracula?,6
post,4pxlu4,2qh72,jokes,false,1466945089,https://old.reddit.com/r/Jokes/comments/4pxlu4/what_is_donald_trumps_biggest_fear/,self.jokes,,Mexican ghosts who can walk through walls.,What is Donald Trump's biggest fear?,5
post,4pxlgs,2qh72,jokes,false,1466944906,https://old.reddit.com/r/Jokes/comments/4pxlgs/the_eu_now_has_1gb_of_free_space/,self.jokes,,#copied,The EU now has 1GB of free space.,5
post,4pxlcd,2qh72,jokes,false,1466944836,https://old.reddit.com/r/Jokes/comments/4pxlcd/why_do_girls_wear_fishnet/,self.jokes,,To show that they're a reel catch.,Why do girls wear fishnet?,1
post,4pxl94,2qh72,jokes,false,1466944797,https://old.reddit.com/r/Jokes/comments/4pxl94/a_man_goes_for_his_first_prostate_exam/,self.jokes,,"""I am sorry doctor, but where can I leave my pants?""

""Right there where I left mine"" - the doctor says",A man goes for his first prostate exam,65
post,4pxkl6,2qh72,jokes,false,1466944459,https://old.reddit.com/r/Jokes/comments/4pxkl6/a_man_went_to_a_meeting_for_premature_ejaculators/,self.jokes,,"but when he arrived there was no one there, he'd come too early. ",A man went to a meeting for premature ejaculators,214
post,4pxk3a,2qh72,jokes,false,1466944213,https://old.reddit.com/r/Jokes/comments/4pxk3a/i_was_gang_raped_by_a_group_of_mimes/,self.jokes,,[removed],I was gang raped by a group of mimes,1
post,4pxk2m,2qh72,jokes,false,1466944199,https://old.reddit.com/r/Jokes/comments/4pxk2m/a_plumber_rings_the_doorbell/,self.jokes,,"""Come in"", says the homeowner, Stacy.

""Hi, I am the plumber, sorry for being a bit late""

""That's fine, my sister must have called for you""

""Alright. So where's that disgusting clogged up mess?""

""Her name actually is Rita, and she's not home at the moment"".",A plumber rings the doorbell,132
post,4pxjfv,2qh72,jokes,false,1466943853,https://old.reddit.com/r/Jokes/comments/4pxjfv/how_do_you_organise_a_space_party/,self.jokes,,You planet.,How do you organise a space party?,7
post,4pxj55,2qh72,jokes,false,1466943683,https://old.reddit.com/r/Jokes/comments/4pxj55/how_do_you_make_a_feminist_mad/,self.jokes,,That isn't funny!,How do you make a feminist mad?,3
post,4pxj2b,2qh72,jokes,false,1466943644,https://old.reddit.com/r/Jokes/comments/4pxj2b/an_indian_girl_is_into_bdsm/,self.jokes,,She's a poppadominatrix,An Indian girl is into BDSM,3
post,4pxix4,2qh72,jokes,false,1466943569,https://old.reddit.com/r/Jokes/comments/4pxix4/donald_trump/,self.jokes,,The joke's in the title.,Donald Trump,0
post,4pxige,2qh72,jokes,false,1466943326,https://old.reddit.com/r/Jokes/comments/4pxige/i_know_a_guy_who_loves_mushrooms/,self.jokes,,...He's a real fun guy!,I know a guy who loves mushrooms..,0
post,4pxiah,2qh72,jokes,false,1466943228,https://old.reddit.com/r/Jokes/comments/4pxiah/what_do_you_call_a_black_priest/,self.jokes,,"holy shit



",What do you call a Black Priest?,0
post,4pxi2z,2qh72,jokes,false,1466943119,https://old.reddit.com/r/Jokes/comments/4pxi2z/friend_left_his_facebook_open_and_his_dad_took/,self.jokes,,[removed],Friend left his Facebook open and his dad took the chance.,1
post,4pxhkr,2qh72,jokes,false,1466942813,https://old.reddit.com/r/Jokes/comments/4pxhkr/why_have_all_remain_voters_suddenly_gotten_so/,self.jokes,,They don't like the taste of being the minority!,Why have all Remain voters suddenly gotten so salty?,0
post,4pxhfb,2qh72,jokes,false,1466942746,https://old.reddit.com/r/Jokes/comments/4pxhfb/what_is_rickon_starks_favourite_band/,self.jokes,,One Direction.,What is Rickon Stark's favourite band ?,5
post,4pxh39,2qh72,jokes,false,1466942561,https://old.reddit.com/r/Jokes/comments/4pxh39/whats_black_and_sits_at_the_top_of_stairs/,self.jokes,,A paraplegic after a house fire.,What's black and sits at the top of stairs?,105
post,4pxh0p,2qh72,jokes,false,1466942529,https://old.reddit.com/r/Jokes/comments/4pxh0p/an_old_man_is_asked_if_he_wears_boxers_or_briefs/,self.jokes,,"He shrugs and says ""Depends.""",An old man is asked if he wears boxers or briefs.,0
post,4pxguf,2qh72,jokes,false,1466942421,https://old.reddit.com/r/Jokes/comments/4pxguf/what_do_you_call_a_dinosaur_that_rapes/,self.jokes,,A sexual predator.,What do you call a dinosaur that rapes?,0
post,4pxgrh,2qh72,jokes,false,1466942368,https://old.reddit.com/r/Jokes/comments/4pxgrh/what_do_you_call_a_dog_in_a_sub/,self.jokes,,"A subwoofer!

Now again: 

What do you call a dog in a sub? 

Chinese food! ",What do you call a dog in a sub?,9
post,4pxg2i,2qh72,jokes,false,1466941956,https://old.reddit.com/r/Jokes/comments/4pxg2i/why_father_cheats_mom/,self.jokes,,Why father cheats mom?,Why father cheats mom?,0
post,4pxfr7,2qh72,jokes,false,1466941773,https://old.reddit.com/r/Jokes/comments/4pxfr7/i_bet_i_can_tell_you_where_you_got_your_shoes/,self.jokes,,You got'em on your feet.,I bet i can tell you where you got your shoes.,26
post,4pxf94,2qh72,jokes,false,1466941482,https://old.reddit.com/r/Jokes/comments/4pxf94/son_dad_what_is_an_idiot/,self.jokes,,[removed],"Son: Dad, what is an idiot?",0
post,4pxf56,2qh72,jokes,false,1466941415,https://old.reddit.com/r/Jokes/comments/4pxf56/whats_the_difference_between_awkward_and_awful/,self.jokes,,"Awkward is finding your mom on Tinder, awful is matching with her",What's the difference between awkward and awful?,29
post,4pxeu6,2qh72,jokes,false,1466941232,https://old.reddit.com/r/Jokes/comments/4pxeu6/why_jews_have_a_big_nose/,self.jokes,,Because the air is free.,Why jews have a big nose?,0
post,4pxekp,2qh72,jokes,false,1466941102,https://old.reddit.com/r/Jokes/comments/4pxekp/whats_the_difference_between_santa_claus_and_a_jew/,self.jokes,,Santa Claus comes DOWN the chimney...,What's the difference between Santa Claus and a jew?,0
post,4pxdhj,2qh72,jokes,false,1466940478,https://old.reddit.com/r/Jokes/comments/4pxdhj/how_do_asians_execute_white_people/,self.jokes,,They cut off their heads using a Gweilotine.,How do Asians execute white people?,0
post,4pxcfk,2qh72,jokes,false,1466939873,https://old.reddit.com/r/Jokes/comments/4pxcfk/i_put_the_sexy_in_dyslexia/,self.jokes,,[removed],I put the sexy in dyslexia.,1
post,4pxcdn,2qh72,jokes,false,1466939842,https://old.reddit.com/r/Jokes/comments/4pxcdn/my_circus_career/,self.jokes,,"My mom and my dad want to send me to a circus to learn how to ride a unicycle(here comes dai boi oh shit waddup)and others so after  a while i got bored and i want to learn sword swallowing so i ask my mom to let me learn sword swallowing and she was so angry and tell me to not talk to her again so i got upset and tell my father,My father laugh at me saying your mother taught you were gay 










do you get it if you dont it is sword swallowing can be related to cock sucking",My Circus career,0
post,4pxc7p,2qh72,jokes,false,1466939739,https://old.reddit.com/r/Jokes/comments/4pxc7p/how_are_white_people_executed_in_asian_countries/,self.jokes,,[deleted],How are white people executed in Asian countries?,1
post,4pxc7a,2qh72,jokes,false,1466939725,https://old.reddit.com/r/Jokes/comments/4pxc7a/what_do_two_bigots_say_to_each_other/,self.jokes,,[removed],What do two bigots say to each other?,1
post,4pxbkj,2qh72,jokes,false,1466939331,https://old.reddit.com/r/Jokes/comments/4pxbkj/what_did_the_feminist_say_when_someone_talked/,self.jokes,,YOUR CHRONO TRIGGERER ME...FUCK YOU THIS IS A FUNNY JOKEFUCKYOUIJUSTWANTYOUTOLOVEMEFUCKYOU,What did the feminist say when someone talked shit about their favorite SNES game?,0
post,4pxbim,2qh72,jokes,false,1466939299,https://old.reddit.com/r/Jokes/comments/4pxbim/a_funny_original_joke_i_came_up_with/,self.jokes,,"Whoops, wrong sub.","A funny, original joke I came up with...",0
post,4pxb9s,2qh72,jokes,false,1466939143,https://old.reddit.com/r/Jokes/comments/4pxb9s/brexit/,self.jokes,,"There is a new slimming product in town. 

It is called Brexit. It'll help you lose a lot of pounds.",Brexit,9
post,4pxaxq,2qh72,jokes,false,1466938929,https://old.reddit.com/r/Jokes/comments/4pxaxq/a_man_was_in_a_state_of_emergency/,self.jokes,,[deleted],A man was in a state of emergency,4
post,4pxaob,2qh72,jokes,false,1466938770,https://old.reddit.com/r/Jokes/comments/4pxaob/a_blind_man_walks_into_a_lesbian_bar/,self.jokes,,"So a blind older gentleman stumbles into a all lesbian bar. They see he is older and blind so they let him stay and have a few drinks. The blind man ask's the bartender ""You want to hear a blonde joke?"" The bartender replies "" Well, I am a blonde, the woman on your right is a defence instructor and she is blonde, and the two woman behind you are marines and they are blonde. Do you still want to tell your joke?"" The blind man responds ""Well not if I have to explain it four times""",A blind man walks into a lesbian bar.,349
post,4pxaj2,2qh72,jokes,false,1466938677,https://old.reddit.com/r/Jokes/comments/4pxaj2/my_lesbian_neighbors_gave_me_a_rolex_for_my/,self.jokes,,"It was mighty kind of them,  but they misunderstood when I said ""I wanna watch""",My lesbian neighbors gave me a Rolex for my birthday,201
post,4px9vr,2qh72,jokes,false,1466938290,https://old.reddit.com/r/Jokes/comments/4px9vr/if_two_atheist_disagreed_whos_wrong/,self.jokes,,[removed],"If two atheist disagreed, who's wrong?",1
post,4px8ih,2qh72,jokes,false,1466937461,https://old.reddit.com/r/Jokes/comments/4px8ih/if_you_ever_get_cold/,self.jokes,,Just stand in a corner. They're usually around 90 degrees!,If you ever get cold...,58
post,4px8dh,2qh72,jokes,false,1466937370,https://old.reddit.com/r/Jokes/comments/4px8dh/michael_jackson/,self.jokes,,I was in Tescos the other day when I saw some bloke who reminded me of Michael Jackson. He came up to me and said 'Never forget Michael Jackson'.,Michael Jackson,1
post,4px7zm,2qh72,jokes,false,1466937116,https://old.reddit.com/r/Jokes/comments/4px7zm/i_married_a_jewish_girl/,self.jokes,,It was the best career move I ever made.,I married a Jewish girl...,4
post,4px7wy,2qh72,jokes,false,1466937070,https://old.reddit.com/r/Jokes/comments/4px7wy/what_is_rickon_starks_favourite_band/,self.jokes,,One Direction,What is Rickon Stark's favourite band?,0
post,4px6yc,2qh72,jokes,false,1466936420,https://old.reddit.com/r/Jokes/comments/4px6yc/what_question_will_get_you_to_the_front_page/,self.jokes,,[removed],What question will get you to the front page?,1
post,4px6fv,2qh72,jokes,false,1466936087,https://old.reddit.com/r/Jokes/comments/4px6fv/ive_been_looking_for_my_exgirlfriends_killer_for/,self.jokes,,[deleted],I've been looking for my ex-girlfriend's killer for past two years,1
post,4px6cc,2qh72,jokes,false,1466936017,https://old.reddit.com/r/Jokes/comments/4px6cc/a_couple_wants_to_have_sex_but_their_son_is_in/,self.jokes,,"The only way to pull off a Sunday afternoon ""quickie "" with their 8-year-old son in the apartment was to send him out on the balcony with a Popsicle and tell him to report on all the neighborhood activities...

""There's a car being towed from the parking lot,"" he shouted.He began his commentary as his parents put their plan into operation.

""An ambulance just drove by!""

""Looks like the Andersons have company,"" he called out.

""Matt's riding a new bike!""

""Looks like the Sanders are moving!""

""Jason is on his skate board!""

After a few moments he announced... ""The Coopers are having sex. Startled, his mother and dad shot up in bed.

Dad cautiously called out...""How do you know they're having sex?"" ""Jimmy Cooper is standing on his balcony with a Popsicle.""
",A couple wants to have sex but their son is in the house.,1113
post,4px65f,2qh72,jokes,false,1466935880,https://old.reddit.com/r/Jokes/comments/4px65f/where_is_macau_located/,self.jokes,,In MaFarm,Where is Macau located?,28
post,4px649,2qh72,jokes,false,1466935855,https://old.reddit.com/r/Jokes/comments/4px649/pigeons/,self.jokes,,"I've just seen a flock of pigeons in army unifoms.

I think it might be a military coo.",Pigeons...,7
post,4px5yo,2qh72,jokes,false,1466935746,https://old.reddit.com/r/Jokes/comments/4px5yo/who_will_pay/,self.jokes,,"If two gays are on a Date for the dinner,Who will pay the bill ?",Who will pay ?,0
post,4px4uz,2qh72,jokes,false,1466935040,https://old.reddit.com/r/Jokes/comments/4px4uz/i_have_a_bad_ping/,self.jokes,,It might be terminal.,I have a bad ping.,6
post,4px4pp,2qh72,jokes,false,1466934939,https://old.reddit.com/r/Jokes/comments/4px4pp/theres_two_fish_in_a_tank_and_one_says/,self.jokes,,"""How do you drive this thing?""","There's two fish in a tank, and one says",7
post,4px4oj,2qh72,jokes,false,1466934917,https://old.reddit.com/r/Jokes/comments/4px4oj/how_are_babies_different_from_feminists/,self.jokes,,Babies grow up and stop crying.,How are babies different from feminists?,14
post,4px4he,2qh72,jokes,false,1466934774,https://old.reddit.com/r/Jokes/comments/4px4he/two_cows_are_scared_of_getting_mad_cow_disease/,self.jokes,,"A cow walks up to another cow and asks 

""Are you scared of Mad Cow Disease?"" 

He replies, shocked

""No, I'm a Duck.""",Two Cows are scared of getting mad cow disease,1
post,4px4gc,2qh72,jokes,false,1466934752,https://old.reddit.com/r/Jokes/comments/4px4gc/who_will_pay/,self.jokes,,[deleted],Who will pay ?,1
post,4px3k7,2qh72,jokes,false,1466934161,https://old.reddit.com/r/Jokes/comments/4px3k7/there_is_a_bomb_going_to_explode_in_321/,self.jokes,,"Holy shit, this blew up! ",There is a bomb going to explode in 3...2...1...,0
post,4px35y,2qh72,jokes,false,1466933940,https://old.reddit.com/r/Jokes/comments/4px35y/ever_since_the_eu_referendum_david_cameron_has/,self.jokes,,People say he's really outgoing,"Ever since the EU referendum, David Cameron has become more friendly than ever..",1
post,4px2xy,2qh72,jokes,false,1466933796,https://old.reddit.com/r/Jokes/comments/4px2xy/my_sister_asked_me_to_take_off_her_clothes/,self.jokes,,[deleted],My sister asked me to take off her clothes.,2
post,4px0km,2qh72,jokes,false,1466932239,https://old.reddit.com/r/Jokes/comments/4px0km/i_have_an_irrational_fear_of_elevators/,self.jokes,,I always feel like they are going to let me down someday.,I have an irrational fear of elevators,12
post,4px0eb,2qh72,jokes,false,1466932142,https://old.reddit.com/r/Jokes/comments/4px0eb/two_mexicans_are_in_a_car_who_drives/,self.jokes,,The police officer,Two mexicans are in a car. Who drives?,32
post,4px0a5,2qh72,jokes,false,1466932063,https://old.reddit.com/r/Jokes/comments/4px0a5/i_wrote_a_book_on_my_sex_change_operation/,self.jokes,,[deleted],I wrote a book on my sex change operation...,1
post,4px02c,2qh72,jokes,false,1466931923,https://old.reddit.com/r/Jokes/comments/4px02c/im_always_suspicious_of_stairs/,self.jokes,,They're usually up to something.,I'm always suspicious of stairs.,12
post,4pwzm1,2qh72,jokes,false,1466931618,https://old.reddit.com/r/Jokes/comments/4pwzm1/3_women_in_a_bar_are_comparing_how_loose_they_are/,self.jokes,,"One claimed they could fit a sausage, another claimed they can fit a cucumber and the other slid down the bar stool. ",3 women in a bar are comparing how loose they are...,120
post,4pwz42,2qh72,jokes,false,1466931299,https://old.reddit.com/r/Jokes/comments/4pwz42/i_asked_a_chinese_girl_for_her_number/,self.jokes,,"I asked a Chinese girl for her number. She replied, ""Sex! Sex! Sex! Free sex tonight!"" I said, ""Wow!"". Then her friend said, ""She means 6663629.""﻿",I asked a Chinese girl for her number,34
post,4pwyp7,2qh72,jokes,false,1466931015,https://old.reddit.com/r/Jokes/comments/4pwyp7/what_do_you_call_a_special_agent_in_a_washing_up/,self.jokes,,Ha bubble 0 7 ,What do you call a special agent in a washing up bottle!?,0
post,4pwyfs,2qh72,jokes,false,1466930850,https://old.reddit.com/r/Jokes/comments/4pwyfs/a_psychic_is_buying_clothes/,self.jokes,,[removed],A psychic is buying clothes.,1
post,4pwyc8,2qh72,jokes,false,1466930788,https://old.reddit.com/r/Jokes/comments/4pwyc8/what_does_a_homeless_man_get_for_christmas/,self.jokes,,[deleted],What does a homeless man get for Christmas?,5
post,4pwyb2,2qh72,jokes,false,1466930768,https://old.reddit.com/r/Jokes/comments/4pwyb2/i_heard_so_many_women_say_its_so_big_i_dont_think/,self.jokes,,But it was mostly on the internet,"I heard so many women say ""it's so big, I don't think it's going to fit"".",0
post,4pwy8e,2qh72,jokes,false,1466930716,https://old.reddit.com/r/Jokes/comments/4pwy8e/what_do_you_call_an_american_communist/,self.jokes,,Manifesto Destiny,What do you call an American communist?,0
post,4pwxy1,2qh72,jokes,false,1466930531,https://old.reddit.com/r/Jokes/comments/4pwxy1/2_inmates_sneer_at_their_new_cellmate/,self.jokes,,"Inmate #1: ""Hey..look at my tattoo. It's a King Cobra. King Cobra! You better watch out, boy.""

The New Inmate says nothing &amp; remains quiet.

Inmate #2: ""Hey..look at my tattoo. It's a Bald Eagle. A Bald Eagle who eats the King Cobra! You better watch out, boy.""

The new inmate slowly gets up &amp; takes of his shirt revealing a large tattoo across his back.

Inmates #1 &amp; #2 look at each other: 
""Oh my god..it's a DRAGON...""

 The new inmate turns around and in a deep &amp; loud voice asks: ""WHAT DID YOU SAY YOUR TATTOOS WERE? HUH!?! TALK!""

Inmate #1: ""Oh..um...err..nothing. just a small, harmless little worm.""

Inmate #2: ""Mm..mine is a cute little chick who eats the cute little worm.""",2 Inmates sneer at their new cellmate..,0
post,4pwxxs,2qh72,jokes,false,1466930528,https://old.reddit.com/r/Jokes/comments/4pwxxs/a_black_man_a_mexican_and_a_chinese_man_all_jump/,self.jokes,,[deleted],"A Black Man, a Mexican, and a Chinese man all jump off a bridge",0
post,4pwxmd,2qh72,jokes,false,1466930325,https://old.reddit.com/r/Jokes/comments/4pwxmd/did_you_hear_those_two_fighting_last_night/,self.jokes,,[deleted],Did you hear those two fighting last night?,0
post,4pwxid,2qh72,jokes,false,1466930258,https://old.reddit.com/r/Jokes/comments/4pwxid/my_girlfriend_like_to_have_anal_sex_4_times_a_day/,self.jokes,,[deleted],My girlfriend like to have anal sex 4 times a day...,0
post,4pwwym,2qh72,jokes,false,1466929953,https://old.reddit.com/r/Jokes/comments/4pwwym/heres_a_nsfw_riddle_i_just_thought_of_while/,self.jokes,,[removed],Here's a NSFW riddle I just thought of while taking a shit.,1
post,4pwwkt,2qh72,jokes,false,1466929736,https://old.reddit.com/r/Jokes/comments/4pwwkt/i_bought_a_llama_on_the_internet_today/,self.jokes,,[deleted],I bought a llama on the internet today,3
post,4pwwf6,2qh72,jokes,false,1466929636,https://old.reddit.com/r/Jokes/comments/4pwwf6/are_you_going_down_there/,self.jokes,,[deleted],Are you going down there?,0
post,4pwwdf,2qh72,jokes,false,1466929609,https://old.reddit.com/r/Jokes/comments/4pwwdf/what_do_you_give_a_girl_who_already_has_everything/,self.jokes,,Antibiotics,What do you give a girl who already has everything?,311
post,4pwvhr,2qh72,jokes,false,1466929007,https://old.reddit.com/r/Jokes/comments/4pwvhr/i_raped_a_blind_woman/,self.jokes,,[deleted],I raped a blind woman...,0
post,4pwvhj,2qh72,jokes,false,1466929002,https://old.reddit.com/r/Jokes/comments/4pwvhj/little_johnny_comes_home_from_school_with_a_note/,self.jokes,,"Johnny's mother reads the note and is astonished as she prepares to scold him.

""Johnny this says you tried to eat Sally, your ant just go around eating people."" She says to the little boy.

Little Johnny looks up at his mother and says ""I know, that's why I got consent first.""",Little Johnny comes home from school with a note.,0
post,4pwvdm,2qh72,jokes,false,1466928934,https://old.reddit.com/r/Jokes/comments/4pwvdm/why_cant_cops_eat_bacon/,self.jokes,,Because that would be cannibalism ,Why can't cops eat bacon?,0
post,4pwv82,2qh72,jokes,false,1466928829,https://old.reddit.com/r/Jokes/comments/4pwv82/every_single_time_i_give_my_heart_to_a_girl/,self.jokes,,She Brexit.,Every single time I give my heart to a girl...,5
post,4pwuzh,2qh72,jokes,false,1466928674,https://old.reddit.com/r/Jokes/comments/4pwuzh/its_time_for_drs_chekup/,self.jokes,,"A man goes to the doctor and says, ""Doctor, wherever I touch, it hurts."" 
The doctor asks, ""What do you mean?"" 
The man says, ""When I touch my shoulder, it really hurts. If I touch my knee - OUCH! When I touch my forehead, it really, really hurts."" 
The doctor says, ""I know what's wrong with you - you've broken your finger!"" ",IT'S TIME FOR DR'S CHEKUP,2
post,4pwuz8,2qh72,jokes,false,1466928671,https://old.reddit.com/r/Jokes/comments/4pwuz8/my_dad_went_to_vietnam/,self.jokes,,"He single-handedly shot and killed 32 north vietnamese. 

Next year we're going on vacation somewhere else.

Edit: spelling",My dad went to Vietnam,3
post,4pwuf5,2qh72,jokes,false,1466928340,https://old.reddit.com/r/Jokes/comments/4pwuf5/why_are_lesbians_bad_cooks/,self.jokes,,because they always eat out...,Why are lesbians bad cooks?,1
post,4pwu2p,2qh72,jokes,false,1466928137,https://old.reddit.com/r/Jokes/comments/4pwu2p/what_was_john_lennons_final_hit/,self.jokes,,The pavement ,What was John Lennons final hit?,5
post,4pwssd,2qh72,jokes,false,1466927335,https://old.reddit.com/r/Jokes/comments/4pwssd/sends_a_remail_to_hillary/,self.jokes,,*Deleted*,*Sends a r/email to Hillary*,0
post,4pwsdv,2qh72,jokes,false,1466927088,https://old.reddit.com/r/Jokes/comments/4pwsdv/hell_isnt_all_that_bad/,self.jokes,,[removed],Hell isn't all that bad!,1
post,4pwr8w,2qh72,jokes,false,1466926443,https://old.reddit.com/r/Jokes/comments/4pwr8w/psychic_buys_clothing/,self.jokes,,"Employee: How about this one?

Psychic: That shirt is too small

Employee: You didn't even try it on

Psychic: I'm a medium",Psychic buys clothing,290
post,4pwq6m,2qh72,jokes,false,1466925817,https://old.reddit.com/r/Jokes/comments/4pwq6m/psychic_buying_clothes/,self.jokes,,[deleted],Psychic Buying Clothes!,1
post,4pwq62,2qh72,jokes,false,1466925810,https://old.reddit.com/r/Jokes/comments/4pwq62/who_makes_the_sandwiches_in_a_lesbian_relationship/,self.jokes,,"Neither, they both eat out.",Who makes the sandwiches in a lesbian relationship?,119
post,4pwo0d,2qh72,jokes,false,1466924525,https://old.reddit.com/r/Jokes/comments/4pwo0d/tifu_i_picked_up_somebody_elses_sandwich_at_subway/,self.jokes,,"Ooops, wrong sub!",[TIFU] I picked up somebody else's sandwich at Subway,16
post,4pwn5l,2qh72,jokes,false,1466924006,https://old.reddit.com/r/Jokes/comments/4pwn5l/do_u_know_whats_a_b_c_d_e_f_g_means/,self.jokes,,[removed],Do u know whats A B C D E F G? means?,1
post,4pwmza,2qh72,jokes,false,1466923904,https://old.reddit.com/r/Jokes/comments/4pwmza/if_10_men_took_2_days_to_build_a_wall_how_long/,self.jokes,,[deleted],"If 10 men took 2 days to build a wall, how long will it take 5 men to build a wall?",0
post,4pwms7,2qh72,jokes,false,1466923803,https://old.reddit.com/r/Jokes/comments/4pwms7/what_do_you_call_a_calculator_with_alcoholics/,self.jokes,,[deleted],What do you call a Calculator with alcoholic's liver disease,1
post,4pwmgi,2qh72,jokes,false,1466923612,https://old.reddit.com/r/Jokes/comments/4pwmgi/if_hillary_is_elected_president/,self.jokes,,[removed],If Hillary is elected president...,0
post,4pwma5,2qh72,jokes,false,1466923518,https://old.reddit.com/r/Jokes/comments/4pwma5/a_train_driver_accidentally_kills_a_man_when_he/,self.jokes,,"Since he killed a person, the court sentences him to death by electrocution chair. For his last meal, he requests a single banana. The prison guard thought it was odd, but gave him the banana, and the man ate it. The next day, the man is strapped onto the electrocution chair and the executioner switches the electricity on. Nothing happened at all. This city has a law that allows a prisoner to walk free if the execution somehow doesn't work, so the train driver was acquitted.

A week later, the train driver miraculously got another job at the train station. However, he drove off the tracks again and killed two people. This man was then arrested immediately and sentenced to death again. For his last meal, the train driver requests two bananas which is fulfilled. The next day, the man is strapped onto the electrocution chair and the executioner turns on the electricity. Nothing happens. So, again, the man is allowed to walk free.

The next week, the train driver somehow managed to get another job at the train station. Again, he drove off the tracks and killed three people. Again, the man was arrested immediately and sentenced to death. This time, for his last meal, the train driver requests three bananas. The exasperated prison guard exclaims, ""Stop! You don't get another banana!"" and takes the train driver to his execution. The train driver once again is strapped onto the chair, and the executioner turns on the electricity. Once again, nothing happens.

The executioner and prison guards are dumbfounded. The train driver laughs and says, ""See? The bananas have nothing to do with my execution— I'm just a bad conductor.""",A train driver accidentally kills a man when he drives off the tracks,65
post,4pwlyo,2qh72,jokes,false,1466923349,https://old.reddit.com/r/Jokes/comments/4pwlyo/hillary_clinton_is_elected_president/,self.jokes,,[removed],Hillary Clinton is elected President.,1
post,4pwltf,2qh72,jokes,false,1466923273,https://old.reddit.com/r/Jokes/comments/4pwltf/anonymous_gets_alzheimers/,self.jokes,,"They sign off: We are Anonymous, we are a legion, we do not forgive, we do not....",Anonymous gets Alzheimer's,0
post,4pwkyp,2qh72,jokes,false,1466922804,https://old.reddit.com/r/Jokes/comments/4pwkyp/why_isnt_infinite_warfare_an_acceptable_password/,self.jokes,,[deleted],"Why isn't ""Infinite Warfare"" an acceptable password?",0
post,4pwkhv,2qh72,jokes,false,1466922572,https://old.reddit.com/r/Jokes/comments/4pwkhv/an_rjokes_mod_an_rconspiracy_mod_an_rnews_mod/,self.jokes,,[deleted],"An r/jokes Mod, an r/conspiracy Mod, &amp; an r/news Mod walk into a bar...",2
post,4pwjnt,2qh72,jokes,false,1466922094,https://old.reddit.com/r/Jokes/comments/4pwjnt/what_do_you_call_a_group_of_senior_japanese/,self.jokes,,Comic Sans,What do you call a group of senior Japanese comedians?,190
post,4pwj0p,2qh72,jokes,false,1466921740,https://old.reddit.com/r/Jokes/comments/4pwj0p/the_ticketmaster_voucher_settlement/,self.jokes,,[removed],The ticketmaster voucher settlement,1
post,4pwiuw,2qh72,jokes,false,1466921662,https://old.reddit.com/r/Jokes/comments/4pwiuw/how_do_you_tell_a_joke_to_a_deaf_person/,self.jokes,,[deleted],How do you tell a joke to a deaf person?,0
post,4pwhla,2qh72,jokes,false,1466921003,https://old.reddit.com/r/Jokes/comments/4pwhla/ive_decided_to_marry_my_midget_girlfriend/,self.jokes,,[deleted],I've decided to marry my midget girlfriend...,1
post,4pwfri,2qh72,jokes,false,1466919992,https://old.reddit.com/r/Jokes/comments/4pwfri/my_mom_just_told_me_she_doesnt_have_a_favorite_kid/,self.jokes,,[deleted],My mom just told me she doesn't have a favorite kid...,3
post,4pwfoq,2qh72,jokes,false,1466919948,https://old.reddit.com/r/Jokes/comments/4pwfoq/did_you_hear_about_the_fish_that_went_deaf/,self.jokes,,"It had to buy a herring aid
",Did you hear about the fish that went deaf?,4
post,4pwfad,2qh72,jokes,false,1466919760,https://old.reddit.com/r/Jokes/comments/4pwfad/yo_mamas_so_fat_she_couldnt_cross_the_road_in_time/,self.jokes,,"...so she went to the ""other side"".","Yo mama's so fat, she couldn't cross the road in time...",0
post,4pwf5v,2qh72,jokes,false,1466919697,https://old.reddit.com/r/Jokes/comments/4pwf5v/my_coworker_sent_me_an_email_about_an_assignment/,self.jokes,,[deleted],My co-worker sent me an email about an assignment.,0
post,4pwev6,2qh72,jokes,false,1466919548,https://old.reddit.com/r/Jokes/comments/4pwev6/why_dont_pc_gamers_get_laid/,self.jokes,,[deleted],Why don't pc gamers get laid,2
post,4pwep1,2qh72,jokes,false,1466919473,https://old.reddit.com/r/Jokes/comments/4pwep1/a_cowboys_vocation/,self.jokes,,"An old cowboy sat down at the bar and ordered a drink. As he sat sipping his drink, a young woman sat down next to him. She turned to the cowboy and asked, ""Are you a real cowboy?""

He replied, ""Well, I've spent my whole life, breaking colts, working cows, going to rodeos, fixing fences, pulling calves, bailing hay, doctoring calves, cleaning my barn, fixing flats, working on tractors, and feeding my dogs, so I guess I am a cowboy.""

She said, ""I'm a lesbian. I spend my whole day thinking about women. As soon as I get up in the morning, I think about women. When I shower, I think about women. When I watch TV, I think about women. I even think about women when I eat. It seems that everything makes me think of women.""

The two sat sipping in silence.

A little while later, a man sat down on the other side of the old cowboy and asked, ""Are you a real cowboy?""

He replied, ""I always thought I was, but I just found out I'm a lesbian.""",A cowboy's vocation,13
post,4pweid,2qh72,jokes,false,1466919377,https://old.reddit.com/r/Jokes/comments/4pweid/can_i_borrow_the_car/,self.jokes,,"There's a family in Alabama that consists of a dad and his son and daughter. One day the daughter goes downstairs to her dad and asks, ""daddy, can I borrow the car tonight to go to my friends party?"" 

The dad replies with ""you know what you've gotta do if you want to borrow the car"" and winked at her.

""But I just sucked your dick last week dad! Please can I just go?"" she retorted. 

Dad says ""you know what ya gotta do hun"" and continues watching his show. 

The daughter thinks about it for a while and decides she really didn't want to miss her friends party. She asks her dad if the offer still stands to which he answered by undoing his belt. 

She reluctantly gets on her knees and goes to start when she looks up and says, ""dad, why does your dick smell like poop?""

Dad replies with ""Oh that's right! Your brother has the car!""",Can I borrow the car?,1
post,4pwdge,2qh72,jokes,false,1466918870,https://old.reddit.com/r/Jokes/comments/4pwdge/why_was_the_tree_in_prison/,self.jokes,,Because it broke every branch of the law.,Why was the tree in prison?,0
post,4pwdgb,2qh72,jokes,false,1466918869,https://old.reddit.com/r/Jokes/comments/4pwdgb/two_beans_on_the_east_coast_of_australia/,self.jokes,,Ended up in Cairns.,Two beans on the east coast of Australia,3
post,4pwd77,2qh72,jokes,false,1466918744,https://old.reddit.com/r/Jokes/comments/4pwd77/what_is_a_terrorist_favorite_pokemon_move/,self.jokes,,Self-Destruct,What is a terrorist favorite Pokemon move?,0
post,4pwchu,2qh72,jokes,false,1466918378,https://old.reddit.com/r/Jokes/comments/4pwchu/what_has_four_wheels_and_flies/,self.jokes,,A Garbage Truck.,"What has four wheels, and flies?",27
post,4pwc3z,2qh72,jokes,false,1466918184,https://old.reddit.com/r/Jokes/comments/4pwc3z/two_priest_walk_into_bar_and_disappointed/,self.jokes,,there are no young boys there.,Two priest walk into bar and disappointed...,0
post,4pwbyv,2qh72,jokes,false,1466918109,https://old.reddit.com/r/Jokes/comments/4pwbyv/what_do_you_call_a_black_pirate/,self.jokes,,[removed],What do you call a black pirate?,0
post,4pwb3j,2qh72,jokes,false,1466917711,https://old.reddit.com/r/Jokes/comments/4pwb3j/a_guy_goes_to_the_doctor_with_a_sore_leg/,self.jokes,,"The doctor runs the normal tests and takes some x-rays. Unable to find the problem he finally decides to listen to the leg with his stethoscope, at the knee he hears ""hey give me $5"" at the calf he hears ""hey give me $10"" at the ankle he hears ""hey give me$15"". He takes off the stethoscope, looks up the patient and says "" I have some bad news, your leg is broke in three places""",A guy goes to the doctor with a sore leg....,75
post,4pw9fy,2qh72,jokes,false,1466916908,https://old.reddit.com/r/Jokes/comments/4pw9fy/adele_is_going_to_have_her_own_childrens_tv_show/,self.jokes,,[deleted],Adele is going to have her own children's tv show...,0
post,4pw9e2,2qh72,jokes,false,1466916887,https://old.reddit.com/r/Jokes/comments/4pw9e2/how_do_you_tell_the_difference_between_a_radical/,self.jokes,,[removed],How do you tell the difference between a radical muslim,0
post,4pw8ma,2qh72,jokes,false,1466916504,https://old.reddit.com/r/Jokes/comments/4pw8ma/started_a_new_religion/,self.jokes,,"Doesn't matter, had sects. ",Started a new religion,10
post,4pw8kf,2qh72,jokes,false,1466916471,https://old.reddit.com/r/Jokes/comments/4pw8kf/hillary_clinton_is_elected_president/,self.jokes,,[removed],Hillary Clinton is elected president,1
post,4pw817,2qh72,jokes,false,1466916202,https://old.reddit.com/r/Jokes/comments/4pw817/so_im_confused_on_where_i_stand_on_masturbation/,self.jokes,,[deleted],So.. I'm confused on where I stand on Masturbation...,0
post,4pw7wp,2qh72,jokes,false,1466916149,https://old.reddit.com/r/Jokes/comments/4pw7wp/what_do_you_call_a_penis_inside_a_potato/,self.jokes,,A dictator,What do you call a Penis inside a Potato?,24
post,4pw7q2,2qh72,jokes,false,1466916057,https://old.reddit.com/r/Jokes/comments/4pw7q2/my_poodle_has_an_amazing_talent_to_whistle_whats/,self.jokes,,"But sadly, you can't hear a dog whistle.",My poodle has an amazing talent to whistle what's on TV/the radio!,0
post,4pw7lj,2qh72,jokes,false,1466916003,https://old.reddit.com/r/Jokes/comments/4pw7lj/somethings_up/,self.jokes,,Has anyone ever seen Donald Trump's and Boris Johnson's hair in the same place at the same time?,Something's up,0
post,4pw79y,2qh72,jokes,false,1466915865,https://old.reddit.com/r/Jokes/comments/4pw79y/you_know_how_i_know_we_are_gonna_have_sex/,self.jokes,,I'm stronger than you!,You know how I know we are gonna have sex?,0
post,4pw6vm,2qh72,jokes,false,1466915679,https://old.reddit.com/r/Jokes/comments/4pw6vm/batman_do_you_bleed/,self.jokes,,"Wonderwoman : No

Batman : ugh.. You forgot to take the pill again didn't you?? ",Batman : Do you bleed??,0
post,4pw3hv,2qh72,jokes,false,1466914056,https://old.reddit.com/r/Jokes/comments/4pw3hv/a_muslim_walks_into_a_gay_bar/,self.jokes,,[removed],A Muslim walks into a gay bar...,1
post,4pw3ba,2qh72,jokes,false,1466913974,https://old.reddit.com/r/Jokes/comments/4pw3ba/two_clowns_walking_in_the_street/,self.jokes,,"The first clown tells the second clown ""Look out, a hole!"".

The seconds responds ""Which hooooooooooooooooooo....""",Two clowns walking in the street,0
post,4pw34z,2qh72,jokes,false,1466913902,https://old.reddit.com/r/Jokes/comments/4pw34z/i_was_at_a_hat_shop_and_the_sign_read_all_caps/,self.jokes,,...and I thought what hypocrites!,"I was at a hat shop and the sign read, ""ALL CAPS MUST GO!""",1
post,4pw2h8,2qh72,jokes,false,1466913616,https://old.reddit.com/r/Jokes/comments/4pw2h8/an_inspector_knocks_on_the_door/,self.jokes,,[removed],an inspector knocks on the door..,2
post,4pw16v,2qh72,jokes,false,1466913009,https://old.reddit.com/r/Jokes/comments/4pw16v/an_inspector_knocks_on_the_door/,self.jokes,,"an inspector knocked on the door.
the six year old boy opened the door and the inspector asked the kid wheres his parents be at? the kid went to the kitchen to call his mom. the mom was cutting a turkey and she accidentally cut her finger. she yells out ""FUCK!"" the six year old asks what does that mean. the mom says ""uh, um it means im cutting a turkey."" the six year old boy then went to go call his dad. the dad was taking a big heavy box to the attic and dropped it on his foot. he screams out ""SHIT"" the six year old boy says what does that mean? the dad says ""it means im taking a box to the attic"" The six year old boy goes back to the inspector and tells the inspector that his mom is fucking a turkey and his dad is taking a shit in the attic. ",an inspector knocks on the door...,0
post,4pw16j,2qh72,jokes,false,1466913004,https://old.reddit.com/r/Jokes/comments/4pw16j/i_hung_out_with_two_guys_named_walter_and_jesse/,self.jokes,,[deleted],I hung out with two guys named Walter and Jesse the other day...,0
post,4pw09w,2qh72,jokes,false,1466912615,https://old.reddit.com/r/Jokes/comments/4pw09w/my_entire_life_is_just_a_test/,self.jokes,,To see whether I'll commit suicide or homicide first.,My entire life is just a test,0
post,4pw08g,2qh72,jokes,false,1466912604,https://old.reddit.com/r/Jokes/comments/4pw08g/inspired_by_chia_pets_a_man_invents_slippers_that/,self.jokes,,[deleted],"Inspired by Chia Pets, a man invents slippers that grow in a similar way. One day he wears them to the store, when a teen comes up to him.",0
post,4pw057,2qh72,jokes,false,1466912563,https://old.reddit.com/r/Jokes/comments/4pw057/chicken/,self.jokes,,[removed],Chicken...,0
post,4pw00h,2qh72,jokes,false,1466912514,https://old.reddit.com/r/Jokes/comments/4pw00h/how_many_mexicans_does_it_take_to_screw_in_a/,self.jokes,,Just Juan.   ,How many Mexicans does it take to screw in a lightbulb?,0
post,4pvzh0,2qh72,jokes,false,1466912284,https://old.reddit.com/r/Jokes/comments/4pvzh0/masturbation_causes_blindness/,self.jokes,,"So one day, my Dad sits me down and tells me ""Son, masturbation is bad and will cause you to go blind. "" 

I had to tell him I was on the other side of the room. ",Masturbation Causes Blindness,0
post,4pvyh1,2qh72,jokes,false,1466911852,https://old.reddit.com/r/Jokes/comments/4pvyh1/those_funny_british/,self.jokes,,[removed],Those Funny British,1
post,4pvyah,2qh72,jokes,false,1466911770,https://old.reddit.com/r/Jokes/comments/4pvyah/jane/,self.jokes,,[removed],Jane...,1
post,4pvxyg,2qh72,jokes,false,1466911629,https://old.reddit.com/r/Jokes/comments/4pvxyg/british_english_will_have_only_3_vowels_now_a_i_o/,self.jokes,,They left E U,British English will have only 3 vowels now A I O,85
post,4pvwv8,2qh72,jokes,false,1466911160,https://old.reddit.com/r/Jokes/comments/4pvwv8/what_do_you_do_when_two_lesbians_make_out_in/,self.jokes,,You get off.,What do you do when two lesbians make out in front of you in a bus?,28
post,4pvv0d,2qh72,jokes,false,1466910336,https://old.reddit.com/r/Jokes/comments/4pvv0d/united_kingdom/,self.jokes,,More like... Divided Kingdom.,United Kingdom,0
post,4pvuhc,2qh72,jokes,false,1466910106,https://old.reddit.com/r/Jokes/comments/4pvuhc/what_do_old_people_with_alzheimers_often_say/,self.jokes,,I don't remember.,What do old people with Alzheimer's often say?,4
post,4pvu95,2qh72,jokes,false,1466910000,https://old.reddit.com/r/Jokes/comments/4pvu95/the_ticket_master_voucher_settlement/,self.jokes,,[removed],The Ticket Master voucher settlement,2
post,4pvtyq,2qh72,jokes,false,1466909862,https://old.reddit.com/r/Jokes/comments/4pvtyq/a_normal_american_guy_bought_the_fastest_and/,self.jokes,," A normal American guy bought the fastest and newest car ever created. He entered the car and turned on the radio; He heard: ""This Is London!"" 
The man said: DAMN this thing is FAST!",A normal American guy bought the fastest and newest car ever created,0
post,4pvssq,2qh72,jokes,false,1466909373,https://old.reddit.com/r/Jokes/comments/4pvssq/why_does_this_certain_race_of_people_drink_so/,self.jokes,,"***""Running in a marathon makes you thirsty....Plus they were all out of the yellow Gatorade!""***

- The race took place in North Dakota....So not a single person was offended, so you shouldn't be either!  ",Why does this certain race of people drink so much of a sugary and grape flavored beverage?,0
post,4pvsip,2qh72,jokes,false,1466909243,https://old.reddit.com/r/Jokes/comments/4pvsip/the_maid_asked_for_a_raise_and_the_wife_was_upset/,self.jokes,,"The maid asked for a raise, and the wife was upset...
She asked, ""Now, Helen, why do you think you deserve a pay increase?""
Helen: ""There are three reasons. The first is that I iron better than you.""
Wife: ""Who said that?""
Helen: ""Your husband.""
Wife: ""Oh.""
Helen: ""The second reason is that I am a better cook than you.""
Wife: ""Who said that?""
Helen: ""Your husband.""
Wife: ""Oh.""
Helen: ""The third reason is that I am better at sex than you.""
Wife: ""Did my husband say that as well?""
Helen: ""No, the gardener did.""
Wife: ""So, how much do you want?""","The maid asked for a raise, and the wife was upset.",2245
post,4pvr1o,2qh72,jokes,false,1466908601,https://old.reddit.com/r/Jokes/comments/4pvr1o/i_was_going_to_make_a_joke_about_brexit/,self.jokes,,But I thought I'd just leave it.,I was going to make a joke about Brexit...,1
post,4pvqug,2qh72,jokes,false,1466908526,https://old.reddit.com/r/Jokes/comments/4pvqug/after_brexit_the_pound_crashed/,self.jokes,,...it's down to ten ounces.,"After #Brexit, the pound crashed...",0
post,4pvq6x,2qh72,jokes,false,1466908252,https://old.reddit.com/r/Jokes/comments/4pvq6x/another_joke_about_drake/,self.jokes,,[deleted],Another joke about Drake,0
post,4pvq6n,2qh72,jokes,false,1466908249,https://old.reddit.com/r/Jokes/comments/4pvq6n/muslim_walks_into_a_night_club_in_florida/,self.jokes,,[removed],Muslim walks into a night club in Florida,0
post,4pvq41,2qh72,jokes,false,1466908218,https://old.reddit.com/r/Jokes/comments/4pvq41/a_man_arrives_to_a_building_answering_to_a_job/,self.jokes,,"A man arrives to a building answering to a job add making nails. 
The boss promptly leads him to the shop which had just a single machine with two levers, two pedals and a rubber pad in the middle. The boss explains: this is the most advanced nail making machine.Pulling the left lever feeds wire to the machine. Pulling the right lever cuts the wire. Stomping the left pedal makes the nail head and stomping the right pedal sharpens the nail tip. Finally you bump the rubber pad with your forehead and it drops the nail into a box. So my friend, I leave you to work. 
The man gets on with the weird dance left hand right hand left foot right foot forehead repeat ... 
About an hour later the boss comes back and asks the man if he's liking his new job to which the man replies ""I like it but I was just thinking..  Maybe you want to stick a broom up my ass so I can start sweeping the shop already, I kind of wanna leave early today"" ",A man arrives to a building answering to a job add making nails. The boss promptly leads him to the shop which had just a single machine,0
post,4pvq0b,2qh72,jokes,false,1466908170,https://old.reddit.com/r/Jokes/comments/4pvq0b/england_may_not_have_a_kidney_bank_but_they_have/,self.jokes,,[removed],"England may not have a kidney bank, but they have a Liverpool.",2
post,4pvpou,2qh72,jokes,false,1466908054,https://old.reddit.com/r/Jokes/comments/4pvpou/a_man_walks_into_a_bar/,self.jokes,,"So a man walks into a local bar. As he walks in he notices a room to the right. This room had four inch plexiglass walls and a faint locking system. In this room it was stacked chest high in 100 dollar bills. He contemplates what it could possibly be for. As he sits down at the bar he asks for a drink. When the bartender pours the drink the man says,         ""Sir, if you don't mind me asking, what is that room for?""                                                                               ""That room contains all the money of the people that failed my bet."" The bartender replies.                  The man continued to drink while wondering what the bet could possibly be. He asked for another drink. This time when the Bartender gets there he asked what the bet was. The bartender simply stated the the bet was for only those brave enough to do the bet, not letting him know what it was. The man was two drinks in and was feeling pretty sure of himself and took the bet.                                       Thus, the bartender told him,""see that man over there in the corner. You have to punch and knock him out with one punch.""                                                 ""I think I can do that. Whiskey,"" said the man.                                  ""But there's more!"" Replied the bartender.                     ""Okay, what else do I have to do? Whiskey!""              ""I have a rabid Pittbull upstairs who needs his teeth pulled out by hand. Also, my 84 year old grand mother is in the room next to it. She has not had an orgasm in 50 years. You need to get her to squirt"".   The man finished another drink, walked right up to nick the brick and knocked him out with one punch. He stumbled upstairs and slammed the door to the dogs room shut. From downstairs all you could hear was growling and whimpering from the dog and the grunting of the man. Then everything went silent. The man started to walk down the stairs again but instead tripped and fell. When he hit the floor, right before he passed out, he looked at the bartender and said,                                                    ""Now where is that old lady who needed her teeth pulled?!""",A man walks into a bar.........,7
post,4pvorr,2qh72,jokes,false,1466907637,https://old.reddit.com/r/Jokes/comments/4pvorr/i_went_to_a_zoo_yesterday_and_the_only_animal_in/,self.jokes,,[deleted],I went to a zoo yesterday and the only animal in the entire zoo was a dog.,0
post,4pvooj,2qh72,jokes,false,1466907604,https://old.reddit.com/r/Jokes/comments/4pvooj/donald_trump_is_elected_president/,self.jokes,,[removed],Donald Trump is elected president,1
post,4pvo13,2qh72,jokes,false,1466907345,https://old.reddit.com/r/Jokes/comments/4pvo13/for_every_upvote_this_gets_my_sheep_and_i_will/,self.jokes,,[deleted],For every upvote this gets my sheep and I will try three thrusts of anal sex.,0
post,4pvnqu,2qh72,jokes,false,1466907221,https://old.reddit.com/r/Jokes/comments/4pvnqu/what_do_you_call_a_sexy_muslim/,self.jokes,,A ji-hottie! ,What do you call a sexy Muslim,34
post,4pvngq,2qh72,jokes,false,1466907097,https://old.reddit.com/r/Jokes/comments/4pvngq/what_do_you_call_a_short_mexican/,self.jokes,,"A paragraph, because they're too short to be an es'e",What do you call a short Mexican?,39
post,4pvmv5,2qh72,jokes,false,1466906838,https://old.reddit.com/r/Jokes/comments/4pvmv5/bernie_sanders_is_elected_president/,self.jokes,,That about covers it.,Bernie Sanders is elected President.,0
post,4pvmf3,2qh72,jokes,false,1466906655,https://old.reddit.com/r/Jokes/comments/4pvmf3/why_do_midgets_laugh_when_they_play_soccer/,self.jokes,,Because the grass tickles their balls.,Why do midgets laugh when they play soccer?,6
post,4pvmae,2qh72,jokes,false,1466906602,https://old.reddit.com/r/Jokes/comments/4pvmae/what_kind_of_bathroom_does_napoleon_use/,self.jokes,,A Waterloo,What kind of bathroom does Napoleon use?,0
post,4pvm0i,2qh72,jokes,false,1466906500,https://old.reddit.com/r/Jokes/comments/4pvm0i/whats_black_white_and_red_and_cant_turn_around_in/,self.jokes,,A nun with a harpoon through her neck,"What's black, white, and red, and can't turn around in a hallway?",0
post,4pvkif,2qh72,jokes,false,1466905867,https://old.reddit.com/r/Jokes/comments/4pvkif/in_every_soap_opera_weve_ever_watched_we_are/,self.jokes,,Didn't stop the Brits from trying,"In every soap opera we've ever watched, we are taught that running away and leaving doesn't solve our problems",3
post,4pvizj,2qh72,jokes,false,1466905194,https://old.reddit.com/r/Jokes/comments/4pvizj/if_two_lesbians_are_on_a_date_who_pays/,self.jokes,,[deleted],"If two lesbians are on a date, who pays?",8223
post,4pvi1z,2qh72,jokes,false,1466904807,https://old.reddit.com/r/Jokes/comments/4pvi1z/every_60_seconds_in_africa/,self.jokes,,a minute passes,Every 60 Seconds in Africa....,3
post,4pvi0i,2qh72,jokes,false,1466904792,https://old.reddit.com/r/Jokes/comments/4pvi0i/a_man_visits_the_doctor_because_of_his_severe/,self.jokes,,"The doctor says, ""It appears that your penis is four inches too long and is pulling on your vocal cords, thereby causing the stutter.""

""D-d-d-oct-t-tor. Wh-ha-a-at c-c-can I d-d-do?""

The doctor tells him that he must remove the extra four inches to relieve the strain.

Six months after the operation, the patient returns for his check-up. ""Doctor, the operation was a success. I no longer stutter, I have a great job and my self-esteem is fantastic. However, my wife says that she misses the great sex we used to have. I was wondering if it is possible to reattach those four inches.""

The doctor hesitates for a minute and then says, ""I d-d-d-on't th-th-think-k-k-k that wo-wo-wo-ould b-be p-p-pos-s-s-ib-b-ble.""
",A man visits the doctor because of his severe stuttering problem.,31
post,4pvhyq,2qh72,jokes,false,1466904771,https://old.reddit.com/r/Jokes/comments/4pvhyq/what_do_you_call_an_optimistic_0/,self.jokes,,A cheery-o!,what do you call an optimistic 0?,9
post,4pvhm2,2qh72,jokes,false,1466904620,https://old.reddit.com/r/Jokes/comments/4pvhm2/does_anyone_have_any_good_tokyo_ghoul_puns/,self.jokes,,I would love if someone would comment some Tokyo Ghoul jokes/puns! Or Attack on Titan... Thx!,Does anyone have any good Tokyo Ghoul puns?,0
post,4pvgt3,2qh72,jokes,false,1466904287,https://old.reddit.com/r/Jokes/comments/4pvgt3/great_britain_has_left_the_eu/,self.jokes,,Now they have a GB of free space,Great Britain has left the EU,1
post,4pvghg,2qh72,jokes,false,1466904165,https://old.reddit.com/r/Jokes/comments/4pvghg/you_have_the_circle_if_light_but_what_do_you_call/,self.jokes,,A noose.,"You have the circle if light, but what do you call the circle of death?",0
post,4pvfz8,2qh72,jokes,false,1466903963,https://old.reddit.com/r/Jokes/comments/4pvfz8/a_guy_called_jim_goes_on_jeopardy_the_round/,self.jokes,,[removed],"A guy called Jim goes on jeopardy, the round begins and the host says...",1
post,4pvfm6,2qh72,jokes,false,1466903801,https://old.reddit.com/r/Jokes/comments/4pvfm6/a_stoner_plumber_walks_into_his_dealers_house/,self.jokes,,"and asks ""where's the shit at?""",A stoner plumber walks into his dealer's house,0
post,4pvete,2qh72,jokes,false,1466903462,https://old.reddit.com/r/Jokes/comments/4pvete/long_visits_to_nature_linked_to_improved_mental/,self.jokes,,Who obviously didn't poll women on Tinder. ,"Long visits to nature linked to improved mental health, study finds. According to new research by Australian and UK environmental scientists.",0
post,4pvdrp,2qh72,jokes,false,1466903045,https://old.reddit.com/r/Jokes/comments/4pvdrp/two_converts_set_off_to_go_join_isis/,self.jokes,,"Hasan and Hussein set off to go join ISIS.  Hasan flew to Istanbul first class, but Hussein was on the no fly list and had to stow away on an empty oil tanker.  But Hasan gifted Hussein a heavy backpack of food and cigarettes to make the trip more bearable.

But when they got to Syria, the ISIS folks found those cigarettes in the backpack and brought them both to a high tower in Raqqa.  

The judge said, ""Hussein, you're pardoned.  But Hasan, we throw you off the tower.""

""But Your Honor,"" Hasan says, ""I'm not even the tobacco junkie!""

""Yeah,"" the judge replies, ""but *he's* on the no fly list.""",Two converts set off to go join ISIS...,3
post,4pvdm7,2qh72,jokes,false,1466902981,https://old.reddit.com/r/Jokes/comments/4pvdm7/usa_is_still_number_one/,self.jokes,,[deleted],U.S.A is still number one..,0
post,4pvc6y,2qh72,jokes,false,1466902385,https://old.reddit.com/r/Jokes/comments/4pvc6y/the_showerhead_and_shower_curtain_are_complaining/,self.jokes,,"Curtain says: I really hate having to just hang here all day.

Showerhead: At least you dont get turned on everytime you see a naked person!",The showerhead and shower curtain are complaining.,6
post,4pvc4d,2qh72,jokes,false,1466902353,https://old.reddit.com/r/Jokes/comments/4pvc4d/i_can_never_talk_to_my_dad_at_breakfast_because/,self.jokes,,I guess you could say he's behind The Times.,I can never talk to my Dad at breakfast because he still reads newspapers.,76
post,4pvbyo,2qh72,jokes,false,1466902273,https://old.reddit.com/r/Jokes/comments/4pvbyo/big_joke/,self.jokes,,[deleted],Big joke !!,0
post,4pvbgh,2qh72,jokes,false,1466902059,https://old.reddit.com/r/Jokes/comments/4pvbgh/whats_the_gayest_dinosaur/,self.jokes,,[deleted],What's the gayest dinosaur?,29
post,4pva8r,2qh72,jokes,false,1466901566,https://old.reddit.com/r/Jokes/comments/4pva8r/death_of_a_general/,self.jokes,,"An army general selected group of personal aids to come along with him when he was visiting a battlefield. At the debriefing, he instructed them that they must follow his instructions no matter what – even if the directions seemed dangerous or counterintuitive. The aids were armed with standard gear and weapons, and they departed for the battlefield. 


Once they arrived, the general decided he wanted to snap a surprise picture of the group with his new camera. He stood up from behind a sandbag, waved his hands, and yelled “Over here! Grin, aids!” 
",Death of a General,3
post,4pva2j,2qh72,jokes,false,1466901503,https://old.reddit.com/r/Jokes/comments/4pva2j/a_good_joke_for_the_engineers_out_there/,self.jokes,,Free time,A good joke for the engineers out there,12
post,4pv9m3,2qh72,jokes,false,1466901321,https://old.reddit.com/r/Jokes/comments/4pv9m3/why_didnt_the_toilet_paper_cross_the_road/,self.jokes,,Because it got stuck in a crack,why didn't the toilet paper cross the road?,3
post,4pv8qv,2qh72,jokes,false,1466900986,https://old.reddit.com/r/Jokes/comments/4pv8qv/real_gutbuster/,self.jokes,,"A woman noticed her husband standing on the bathroom scale, sucking in his stomach. “Ha­­! That’s not going to help,” she said.

“Sure, it does,” he said. “It’s the only way I can see the numbers.”

",real gut-buster,3
post,4pv8mf,2qh72,jokes,false,1466900936,https://old.reddit.com/r/Jokes/comments/4pv8mf/long_death_of_a_general/,self.jokes,,[deleted],[long] Death of a General,1
post,4pv8hh,2qh72,jokes,false,1466900890,https://old.reddit.com/r/Jokes/comments/4pv8hh/some_notes_for_the_mods/,self.jokes,,[removed],Some notes for the mods,1
post,4pv8f0,2qh72,jokes,false,1466900864,https://old.reddit.com/r/Jokes/comments/4pv8f0/a_buddhist_monk_walks_up_to_a_hot_dog_stand_and/,self.jokes,,"""Make me one with everything""",A Buddhist monk walks up to a hot dog stand and says,1
post,4pv7ci,2qh72,jokes,false,1466900415,https://old.reddit.com/r/Jokes/comments/4pv7ci/the_grass_is_always_greener_on_the_other_side/,self.jokes,,[deleted],The grass is always greener on the other side..,0
post,4pv6wq,2qh72,jokes,false,1466900233,https://old.reddit.com/r/Jokes/comments/4pv6wq/her_knickers_come_down_faster_than_the_pound_on/,self.jokes,,[removed],Her knickers come down faster than the pound on Brexit night.,1
post,4pv6tp,2qh72,jokes,false,1466900199,https://old.reddit.com/r/Jokes/comments/4pv6tp/did_you_hear_about_the_two_men_who_were_arrested/,self.jokes,,They each got six months,Did you hear about the two men who were arrested for stealing a calendar?,14
post,4pv6mf,2qh72,jokes,false,1466900111,https://old.reddit.com/r/Jokes/comments/4pv6mf/a_man_walks_into_a_bar/,self.jokes,,Ouch!,A man walks into a bar,9
post,4pv69r,2qh72,jokes,false,1466899969,https://old.reddit.com/r/Jokes/comments/4pv69r/you_might_be_a_redneck_if/,self.jokes,,"The ufo hotline limits you to 1 call per day,
You mow your yard and find a car,
Have less teeth than your 2 year old,
Walk your child to school because your in the same grade,
See a sign saying ""say no to crack"" and you pull your pants,
Your dog and wallet are both on a chain,
People ask to hunt in your yard,
Someone shows up to your house once a day mistakenly thinking your having a yard sale.",You might be a redneck if...,0
post,4pv66y,2qh72,jokes,false,1466899934,https://old.reddit.com/r/Jokes/comments/4pv66y/there_is_a_spice_shortage/,self.jokes,,"There is a shortage of spices all around the world. One entrepreneur saw the shortage coming and stocked up. His advisor was pushing to sell it soon so that people could have all of their favorite dishes. The entrepreneur looked at his advisor and said ""what's the rush? We've got all the thyme in the world.""",There is a spice shortage...,61
post,4pv5v2,2qh72,jokes,false,1466899816,https://old.reddit.com/r/Jokes/comments/4pv5v2/what_do_you_call_a_potato_in_a_polling_room/,self.jokes,,[removed],what do you call a potato in a polling room?,1
post,4pv5p6,2qh72,jokes,false,1466899749,https://old.reddit.com/r/Jokes/comments/4pv5p6/two_guys_are_playing_guess_what/,self.jokes,,[deleted],"Two guys are playing ""Guess what""",0
post,4pv5h7,2qh72,jokes,false,1466899654,https://old.reddit.com/r/Jokes/comments/4pv5h7/mr_and_mrs_needle_were_so_proud_of_their_son_when/,self.jokes,,"While growing up, he was a little prick.",Mr. and Mrs. Needle were so proud of their son when he grew up to be an upstanding citizen.,0
post,4pv50s,2qh72,jokes,false,1466899478,https://old.reddit.com/r/Jokes/comments/4pv50s/i_like_my_women_like_i_like_my_coffee/,self.jokes,,tied up in burlap and thrown over the back of a donkey.,"I like my women like I like my coffee,",0
post,4pv4hb,2qh72,jokes,false,1466899263,https://old.reddit.com/r/Jokes/comments/4pv4hb/i_took_a_shower_today/,self.jokes,,[deleted],I took a shower today.,0
post,4pv46e,2qh72,jokes,false,1466899145,https://old.reddit.com/r/Jokes/comments/4pv46e/whats_the_difference_between_a_hooker_and_a_drug/,self.jokes,,A hooker can wash her crack and sell it again.,What's the difference between a hooker and a drug dealer?,0
post,4pv3cs,2qh72,jokes,false,1466898805,https://old.reddit.com/r/Jokes/comments/4pv3cs/a_few_puns/,self.jokes,,"Q.Why was the toilet paper rolling down the mountain?
A.To get to the bottom!

I heard Apple is designing a new automatic car. But they're having trouble installing windows.

What did the sea say to the sand? Nothing, it simply waved.

I never knew eggs were good for the eyes, but my cousin claims they gave him eggcelent vision.



",A Few Puns,3
post,4pv3bo,2qh72,jokes,false,1466898791,https://old.reddit.com/r/Jokes/comments/4pv3bo/what_do_you_call_an_army_of_toddlers/,self.jokes,,Infantry. ,What do you call an army of toddlers?,34
post,4pv242,2qh72,jokes,false,1466898291,https://old.reddit.com/r/Jokes/comments/4pv242/how_can_you_tell_if_someone_is_from_texas/,self.jokes,,[deleted],How can you tell if someone is from Texas?,1
post,4pv0v6,2qh72,jokes,false,1466897757,https://old.reddit.com/r/Jokes/comments/4pv0v6/i_like_my_comedic_timing_like_my_pizza_delivery/,self.jokes,,With pepperoni.,I like my comedic timing like my pizza delivery,0
post,4pv0px,2qh72,jokes,false,1466897705,https://old.reddit.com/r/Jokes/comments/4pv0px/what_do_you_call_a_wookiee_banker/,self.jokes,,[deleted],What do you call a wookiee banker?,1
post,4puzws,2qh72,jokes,false,1466897394,https://old.reddit.com/r/Jokes/comments/4puzws/three_guys_on_a_corner_when_a_cop_pulls_up/,self.jokes,,[deleted],Three guys on a corner when a cop pulls up,2
post,4puzuo,2qh72,jokes,false,1466897367,https://old.reddit.com/r/Jokes/comments/4puzuo/what_was_bruce_lees_favorite_drink/,self.jokes,,Waattaaah!,What was Bruce Lee's favorite drink?,9
post,4puze3,2qh72,jokes,false,1466897157,https://old.reddit.com/r/Jokes/comments/4puze3/was_in_tesco_this_morning_when_the_cashier_asked/,self.jokes,,[deleted],"Was in tesco this morning, when the cashier asked the foreign couple in front of me if they needed help packing their bags.",3
post,4puz5u,2qh72,jokes,false,1466897047,https://old.reddit.com/r/Jokes/comments/4puz5u/my_grandpa_told_me_this_one/,self.jokes,,"So an older couple is discussing the inevitable matter of death. The wife asks her husband, ""If I die before you do, will you remarry?"" To which the husband replies, ""Well, I don't want to be lonely for the rest of my life, so yes."" The wife then asks, ""What about the house? Will you live in the same house?"" And the husband says, ""Well, I suppose, I mean, it's already paid for."" The wife, getting a little protective, asks, ""And what about my car? Will she drive my car?"" The husband says again, ""Well, it's already paid for..."" The wife, annoyed at this point, shoots, ""What about my golf clubs?!?"" And the husband says, ""Oh, no. She's left handed.""",My grandpa told me this one...,77
post,4puyx5,2qh72,jokes,false,1466896943,https://old.reddit.com/r/Jokes/comments/4puyx5/koale_who_smokes_weed/,self.jokes,,"Long time ago there was a Koala. Sitting on top of his tree where he's always chilling. But today it's different. He is bored as f*ck. So out of boredom he rolled a blunt,

After smoking for like 5 minutes, a lizzard shows up passing by the tree. ""Wait, I know that smell. Hey! Watcha doing?"" he said while looking up. ""Smoking some weed because I""m bored man. U wanna join me mate?"" ""Sure!"" said the lizzard as he climbed up and up untill he reached the Koala.

20 minutes has passed. The lizzard said, after he laughed at a joke koala told: ""Damn I'm so thirsthy. Do u have any water?"" ""Sure"" said the koala. ""Just go down, Then go to your right there about the 10th tree on your left. There's a lake with plenty of water."" ""Thanks!"" said the lizzard as he climbed down the tree and searched for the lake.""

He's really enjoying the water as he drank. But then! The unexpected happend. He fell in the water! Unable to swim, he almost drowned. A big crocodile who saw what happend jumped in the water to save the little lizzard. ""DUDE! U know u can't swim, what are u doing here in the water?"" ""I""m so sorry but i was smoking weed with my koala friend, and I got thursty so I went for a drink."" ""Weed?"" asked the aligater. And where is this koala bear? ""Oh he is over there. about 10 trees further then to your left.""

The koala, smoking his last little bit of weed, looks down an sees the crocodile. ""Goddamn, How much water did u drank?""",Koale who smokes weed,15
post,4puyn2,2qh72,jokes,false,1466896834,https://old.reddit.com/r/Jokes/comments/4puyn2/watch_out_for_children_on_the_road/,self.jokes,,They're terrible drivers. ,Watch out for children on the road.,13
post,4puyjt,2qh72,jokes,false,1466896803,https://old.reddit.com/r/Jokes/comments/4puyjt/whats_at_the_end_of_every_movie/,self.jokes,,Insert coin,What's at the end of every movie?,0
post,4puxt0,2qh72,jokes,false,1466896482,https://old.reddit.com/r/Jokes/comments/4puxt0/everybody_type_in_chat_alex_is_a_stupid_nigger/,self.jokes,,[removed],Everybody type in chat Alex is a stupid nigger,1
post,4puxi3,2qh72,jokes,false,1466896360,https://old.reddit.com/r/Jokes/comments/4puxi3/what_do_you_call_a_joke_without_a_punchline/,self.jokes,,[removed],What do you call a joke without a punchline?,1
post,4puxdy,2qh72,jokes,false,1466896316,https://old.reddit.com/r/Jokes/comments/4puxdy/have_you_seen_the_german_comedian_that_tells/,self.jokes,,I hear he's the wurst.,Have you seen the German Comedian that tells nothing but jokes about Sausage?,1
post,4puwl8,2qh72,jokes,false,1466896036,https://old.reddit.com/r/Jokes/comments/4puwl8/i_saw_a_blind_man_walking_down_the_street_one/,self.jokes,,"I saw a blind man walking down the street one morning and as he passes by a fish market, he shouts ""Good morning ladies!!!"" ",I saw a blind man walking down the street one morning...,1
post,4puw8w,2qh72,jokes,false,1466895915,https://old.reddit.com/r/Jokes/comments/4puw8w/what_type_of_hepatitis_do_canadians_the_fonz_get/,self.jokes,,[deleted],What type of hepatitis do Canadians the Fonz get?,1
post,4puvxe,2qh72,jokes,false,1466895798,https://old.reddit.com/r/Jokes/comments/4puvxe/he_was_the_best_astronomer_in_the_world_he_could/,self.jokes,,He was depressed because he never got to explore HER black hole.,"He was the best astronomer in the world, he could even explore black holes, but...",0
post,4puvuq,2qh72,jokes,false,1466895775,https://old.reddit.com/r/Jokes/comments/4puvuq/colonoscopy/,self.jokes,,[deleted],Colonoscopy,6
post,4puvno,2qh72,jokes,false,1466895712,https://old.reddit.com/r/Jokes/comments/4puvno/hillary_clinton_is_elected_president/,self.jokes,,[removed],Hillary Clinton is elected president,1
post,4puvf7,2qh72,jokes,false,1466895627,https://old.reddit.com/r/Jokes/comments/4puvf7/why_did_the_weather_channel_go_out_of_business/,self.jokes,,Let me know your guesses in the comment section below,Why did the Weather channel go out of business?,0
post,4puv6y,2qh72,jokes,false,1466895529,https://old.reddit.com/r/Jokes/comments/4puv6y/youre_a_carrot/,self.jokes,,"I wish, I'd be easier on the eyes.",You're a Carrot,0
post,4puuum,2qh72,jokes,false,1466895393,https://old.reddit.com/r/Jokes/comments/4puuum/get_hitched_or_die_trying/,self.jokes,,[removed],Get hitched or die trying,1
post,4puu3z,2qh72,jokes,false,1466895112,https://old.reddit.com/r/Jokes/comments/4puu3z/trump_is_elected_president/,self.jokes,,[removed],Trump is elected president...,1
post,4putuc,2qh72,jokes,false,1466895008,https://old.reddit.com/r/Jokes/comments/4putuc/women_say_men_are_warm_even_in_winter/,self.jokes,,[deleted],Women say men are warm even in winter.,0
post,4putrh,2qh72,jokes,false,1466894977,https://old.reddit.com/r/Jokes/comments/4putrh/a_carrot_a_pineapple_and_a_melon_walk_into_a_bar/,self.jokes,,"The melon asks the bartender 
 
""can I have a glass of water?"". 

The bartender, scared and confused as to how he is seeing 3 walking and talking fruit and veg, whips out his cock and starts to gently rub it.

""Excuse me sir, that's a mighty large pipe you got yourself!"" Says the Carrot.

""Oh this lil thang?"", the bartender moans, ""my papa showed me how to use it right......mee hoy minoy"".","A carrot, a pineapple and a melon walk into a bar...",0
post,4putnf,2qh72,jokes,false,1466894928,https://old.reddit.com/r/Jokes/comments/4putnf/why_do_asian_women_have_small_boobs/,self.jokes,,[deleted],Why do Asian women have small boobs?,2
post,4puth8,2qh72,jokes,false,1466894862,https://old.reddit.com/r/Jokes/comments/4puth8/this_woman_i_met_last_night_says_she_wants_a_guy/,self.jokes,,Yet when I tapped on the kitchen window uninvited late at night dressed as a clown it is all panic and screaming.,"This woman I met last night says she wants a guy who is ""spontaneous and fun"".",18
post,4pusgo,2qh72,jokes,false,1466894467,https://old.reddit.com/r/Jokes/comments/4pusgo/an_irashman_walks_out_of_a_bar/,self.jokes,https://www.reddit.com/r/Jokes/comments/4pusgo/an_irashman_walks_out_of_a_bar/,,An irashman walks out of a bar...,4
post,4pusam,2qh72,jokes,false,1466894400,https://old.reddit.com/r/Jokes/comments/4pusam/if_you_are_fat/,self.jokes,,"go to the UK, you will lose a couple of pounds ",If you are fat...,0
post,4pus1o,2qh72,jokes,false,1466894306,https://old.reddit.com/r/Jokes/comments/4pus1o/why_do_milking_stools_only_have_three_legs/,self.jokes,,'Cause the cow has the udder,Why do milking stools only have three legs?,15
post,4purxl,2qh72,jokes,false,1466894262,https://old.reddit.com/r/Jokes/comments/4purxl/a_man_and_his_dog_are_sitting_at_home/,self.jokes,,[removed],a Man and his dog are sitting at home...,1
post,4purfl,2qh72,jokes,false,1466894048,https://old.reddit.com/r/Jokes/comments/4purfl/how_do_you_call_a_20_years_old_cat_an_antikitty/,self.jokes,,[removed],How do you call a 20 years old cat ? -An antikitty,1
post,4puqyz,2qh72,jokes,false,1466893849,https://old.reddit.com/r/Jokes/comments/4puqyz/married_10_times_still_a_virgin/,self.jokes,,"A lawyer married a woman who had previously divorced ten husbands. 

On their wedding night, she told her new husband, ""Please be gentle, I'm still a virgin."" 

""What?"" said the puzzled groom. 

""How can that be if you've been married ten times?"" 

""Well, Husband #1 was a sales representative: he kept telling me how great it was going to be. 

Husband #2 was in software services: he was never really sure how it was supposed to function, but he said he'd look into it and get back to me. 

Husband #3 was from field services: he said everything checked out diagnostically but he just couldn't get the system up. 

Husband #4 was in telemarketing: even though he knew he had the order, he didn't know when he would be able to deliver. 

Husband #5 was an engineer: he understood the basic process but wanted three years to research, implement, and design a new state-of-the-art method. 

Husband #6 was from finance and administration: he thought he knew how, but he wasn't sure whether it was his job or not. 

Husband #7 was in marketing: although he had a nice product, he was never sure how to position it. 

Husband #8 was a psychologist: all he ever did was talk about it. 

Husband #9 was a gynecologist: all he did was look at it. 

Husband #10 was a stamp collector: all he ever did was... God! I miss him! But now that I've married you, I'm really excited!"" 

""Good,"" said the new husband, ""but, why?"" 

""You're a lawyer. This time I know I'm gonna get screwed!""","Married 10 times, still a virgin",47
post,4puqkn,2qh72,jokes,false,1466893686,https://old.reddit.com/r/Jokes/comments/4puqkn/dirty_a_man_starts_dating_a_somewhat_butch_woman/,self.jokes,,"She's got a great personality and they hit it off, but he begins to hear rumors about town that she's actually a man.  She's a bit shy, and they have yet to be intimate, so he's not 100% sure of her gender and it begins to bother him a bit.

One night, he takes her on a date to a drive-in movie theater.  As they watch the movie, she begins to squirm in her seat and says ""I've really got to go to the bathroom"".  Thinking quickly, he says ""I saw a sign that says the bathrooms are out of order, so you'll have to go in the bushes.""  She replies ""I don't care, I have to go"" and hops out of the car and disappears into the bushes.

He waits a few seconds, then quietly slips out of the car and creeps towards her, hoping to get a glimpse of whatever equipment she (he?) is packing.  Sure enough, he sees her crouching slightly behind a bush, and spots something long and thin dangling between her legs.

""Ah ha!"" he yells and reflexively grasps the dangling object.  She screams and says, ""You didn't tell me you're a peeping tom!""  He replies queasily, looking at his hand in disgust, ""You didn't tell me you had to take a shit!""","**Dirty** A Man Starts Dating A Somewhat ""Butch"" Woman",19
post,4puq2b,2qh72,jokes,false,1466893497,https://old.reddit.com/r/Jokes/comments/4puq2b/how_do_you_know_when_the_woman_is_lying/,self.jokes,,[deleted],How do you know when the woman is lying?,0
post,4puorq,2qh72,jokes,false,1466892978,https://old.reddit.com/r/Jokes/comments/4puorq/what_day_do_people_eat_on/,self.jokes,,Tuesday,What day do people eat on?,0
post,4puomi,2qh72,jokes,false,1466892920,https://old.reddit.com/r/Jokes/comments/4puomi/im_no_weatherman/,self.jokes,,[deleted],I'm no weatherman...,1
post,4puohy,2qh72,jokes,false,1466892864,https://old.reddit.com/r/Jokes/comments/4puohy/did_you_know_frogs_can_jump_higher_than_houses/,self.jokes,,"This is for two reasons:

1. Frogs have extremely strong hind legs.

2. Houses can't jump.",Did you know frogs can jump higher than houses?,0
post,4puodn,2qh72,jokes,false,1466892815,https://old.reddit.com/r/Jokes/comments/4puodn/a_texan_donald_trump_and_a_new_mexican_are/,self.jokes,,"They all immediately grab for it, and each get a hand on it. 

As they each struggle to take it from the other two, a genie pops out. The genie says, ""You have woken me from my slumber, and I shall give you three wishes. Since you each have a hand on the lamp, you will get one wish a piece.""

The Donald Trump goes first. He says, ""I want all the Mexicans permanently out of the United States and back in Mexico.""

""So it shall be,"" replies the genie, and suddenly every single Mexican is gone from the US and back in Mexico. 

The Texan then shouts, ""I'm next. You're telling me that all the Mexicans are gone from the US?"" ""Yes,"" replies the genie. The Texan replies, ""OK,I want a 500 foot tall wall around the entire state of Texas so nothing can get in or out.""

""So it shall be,"" replies the genie. Suddenly, a wall begins rising from the ground around the borders of Texas, and the Texan yells out with happiness. 

Lastly, it was the New Mexican's turn. He thinks for a moment, and then asks the genie, ""you're saying there is now a 500 foot wall all around Texas and nothing can get in or out?"" ""Yes,"" replies the genie, ""what is your wish?""

The New Mexican then says to the genie with a huge smile, ""fill it with water."" 

.

.

I was in the ""Texit"" thread when I remembered this joke. I updated the characters to fit 2016. :)

Edit to fix typo","A Texan, Donald Trump, and a New Mexican are walking along when they stumble upon a gold lamp...",204
post,4puo4y,2qh72,jokes,false,1466892711,https://old.reddit.com/r/Jokes/comments/4puo4y/whats_worse_than_dropping_your_ice_cream/,self.jokes,,The Holocaust.,What's worse than dropping your ice cream?,0
post,4punap,2qh72,jokes,false,1466892386,https://old.reddit.com/r/Jokes/comments/4punap/would_you_rather_have_parkinsons_or_dementia/,self.jokes,,Parkinson's I'd rather spill half a beer than forget where I put a full one.,Would you rather have Parkinson's or dementia...,0
post,4pumtd,2qh72,jokes,false,1466892193,https://old.reddit.com/r/Jokes/comments/4pumtd/how_do_you_know_youre_in_scotland/,self.jokes,,There's a Chinese restaurant called Bon Appetit,How do you know you're in Scotland?,0
post,4pumkr,2qh72,jokes,false,1466892096,https://old.reddit.com/r/Jokes/comments/4pumkr/how_do_you_know_when_the_woman_is_lying_to_you/,self.jokes,,[deleted],How do you know when the woman is lying to you?,1
post,4pum11,2qh72,jokes,false,1466891866,https://old.reddit.com/r/Jokes/comments/4pum11/what_came_first_the_chicken_or_the_egg/,self.jokes,,The chicken. Did it 7 times in a row in fact.,What came first? The chicken or the egg?,0
post,4pukrd,2qh72,jokes,false,1466891370,https://old.reddit.com/r/Jokes/comments/4pukrd/tarzan_said_to_george_of_the_jungle/,self.jokes,,"“George, I don’t get it. I’m better at swinging from vines, but you’re still more popular than me. What can I do to be as entertaining as you?”

George shrugged and said, 

“You just have to tree harder.""
",Tarzan said to George of the Jungle,0
post,4puk9k,2qh72,jokes,false,1466891190,https://old.reddit.com/r/Jokes/comments/4puk9k/what_do_you_call_a_male_who_doesnt_know_how_to/,self.jokes,,[deleted],What do you call a male who doesn't know how to use a condom?,37
post,4pujv2,2qh72,jokes,false,1466891038,https://old.reddit.com/r/Jokes/comments/4pujv2/this_probably_counts_as_a_joke_i_certainly/,self.jokes,,[deleted],This probably counts as a joke. I certainly laughed. (Read the whole thing),1
post,4pujtd,2qh72,jokes,false,1466891014,https://old.reddit.com/r/Jokes/comments/4pujtd/i_like_my_girlfriends_like_i_like_my_scotch/,self.jokes,,Twelve years old and mixed up with coke ,I like my girlfriends like I like my scotch,11
post,4pujmq,2qh72,jokes,false,1466890946,https://old.reddit.com/r/Jokes/comments/4pujmq/i_plagiarized_a_book_about_native_americans/,self.jokes,,I eventually got siouxed.,I plagiarized a book about native Americans...,10
post,4pujjt,2qh72,jokes,false,1466890908,https://old.reddit.com/r/Jokes/comments/4pujjt/what_do_you_call_it_when_a_king_gets_a_vasectomy/,self.jokes,,A heir cut,What do you call it when a King gets a vasectomy?,1
post,4pujjb,2qh72,jokes,false,1466890904,https://old.reddit.com/r/Jokes/comments/4pujjb/what_can_destroy_a_great_library_the_fastest/,self.jokes,,A Kindle.,What can destroy a Great Library the fastest?,0
post,4pujdi,2qh72,jokes,false,1466890844,https://old.reddit.com/r/Jokes/comments/4pujdi/whats_the_difference_between_a_porcupine_and_a_bmw/,self.jokes,,A porcupine has pricks on the outside.,Whats the difference between a porcupine and a BMW?,68
post,4puj5u,2qh72,jokes,false,1466890767,https://old.reddit.com/r/Jokes/comments/4puj5u/i_entered_a_pun_contest/,self.jokes,,...on the radio last week.  I won.,I entered a pun contest...,0
post,4puj3z,2qh72,jokes,false,1466890746,https://old.reddit.com/r/Jokes/comments/4puj3z/whats_common_between_reddit_and_a_bad_restaurant/,self.jokes,,"all of our servers are busy right now

please try again in a minute",What's common between Reddit and a bad restaurant?,0
post,4puiwc,2qh72,jokes,false,1466890655,https://old.reddit.com/r/Jokes/comments/4puiwc/british_english/,self.jokes,,"Now British English will have only 3 vowels
**A I O ... **

as it has left E U .... :)",British English,25
post,4puiwb,2qh72,jokes,false,1466890655,https://old.reddit.com/r/Jokes/comments/4puiwb/scientists_have_discovered_that_mothers_are_the/,self.jokes,,"
Because Force = ma.",Scientists have discovered that mothers are the driving force behind their children.,7
post,4puim2,2qh72,jokes,false,1466890533,https://old.reddit.com/r/Jokes/comments/4puim2/_/,self.jokes,,[removed],£,1
post,4puhjn,2qh72,jokes,false,1466890130,https://old.reddit.com/r/Jokes/comments/4puhjn/brexit_joke_for_teh_luls/,self.jokes,,"David cameron was tripping on lsd

""oh my god guys I see a tree""

""come over here tree""

but the tree refused to move.

After some time david cameron decided he would marry the tree

""tree will you marry me?""

but the tree did not respond

David cameron started to get paranoid that the tree would not marry him

""HMM perhaps its time for a brexit""

the tree responded, ""Cameron thats not a good idea, paranoia is not a security, a security is secure, you will fk up the stock market you dingnut""

""Tree I no longer wish to marry you""

And that is the story of brexit",Brexit joke for teh luls,0
post,4puhjb,2qh72,jokes,false,1466890126,https://old.reddit.com/r/Jokes/comments/4puhjb/my_deodorant_is_called_states_evidence/,self.jokes,,Part of the Wetness Protection program.,"My deodorant is called ""state's evidence""...",5
post,4puhbm,2qh72,jokes,false,1466890044,https://old.reddit.com/r/Jokes/comments/4puhbm/i_like_my_woman_like_i_like_my_coffee/,self.jokes,,Ground up and in the freezer,I like my woman like I like my coffee,1
post,4pugvq,2qh72,jokes,false,1466889862,https://old.reddit.com/r/Jokes/comments/4pugvq/if_you_are_fat/,self.jokes,,"If you are far, go to the UK, you will lose a couple of pounds ",If you are fat...,0
post,4pugop,2qh72,jokes,false,1466889770,https://old.reddit.com/r/Jokes/comments/4pugop/who_is_the_pound_for_pound_best_fighter_currently/,self.jokes,,Definitely not the UK ,Who is the pound for pound best fighter currently?,0
post,4pug2w,2qh72,jokes,false,1466889433,https://old.reddit.com/r/Jokes/comments/4pug2w/i_was_so_sad_when_i_heard_gandhi_was_a_racist/,self.jokes,,[deleted],I was so sad when I heard Gandhi was a racist....,6
post,4puf8k,2qh72,jokes,false,1466889125,https://old.reddit.com/r/Jokes/comments/4puf8k/midget/,self.jokes,,[removed],Midget,1
post,4puf7b,2qh72,jokes,false,1466889112,https://old.reddit.com/r/Jokes/comments/4puf7b/three_young_students_finished_a_biology_exam_and/,self.jokes,,"One got an A, the other a B and the third an F. They see a girl walking down the street. The A student says: Gooorrrr I'd love to put my hands on her tits and rub my dick against her ass. The B student says: Gooorrrr I'd love to put my fingers up her panties and finger her. The F student says: Gooorrrr I'd love to pull up her skirt and lick her balls.",Three young students finished a biology exam and are walking down the street.,0
post,4puf59,2qh72,jokes,false,1466889097,https://old.reddit.com/r/Jokes/comments/4puf59/an_85yearold_man_had_to_take_a_sperm_count_for/,self.jokes,,"The doctor gave the man a jar and said, ""Take this jar home and bring back a semen sample tomorrow."" The next day the 85-year-old man reappeared at the doctor's office and gave him the jar, which was as clean and empty as on the previous day. The doctor asked, what happened and the man explained. ""Well, doc, it's like this--first I tried with my right hand, but nothing. Then I tried with my left hand, but still nothing. Then I asked my wife for help. She tried with her right hand, then with her left, still nothing. She tried with her mouth, first with the teeth in, then with her teeth out, still nothing. We even called up Arleen, the lady next door and she tried too, first with both hands, then an armpit, and she even tried squeezin' it between her knees, but still nothing."" The doctor was shocked! ""You asked your neighbor?"" The old man replied, ""Yep, none of us could get the jar open.",An 85-year-old man had to take a sperm count for his physical exam,288
post,4puebo,2qh72,jokes,false,1466888791,https://old.reddit.com/r/Jokes/comments/4puebo/one_day_the_red_and_white_knight_on_a_black_and/,self.jokes,,"A few moments later a guard answered, he looked at the Red and White Knight on a Black and White Horse and said ""This is the castle of the king of England who are you?"".

The Red and White Knight on a Black and White Horse got down off his horse and said ""I am the Red and White Knight on a Black and White Horse, and I want to see the King"" 

The guard looked at him for a while and said ""Red and White Knight on a Black and White Horse, I will ask the king if he will grant you an audience"".

The guard went through the castle and to the kings throne room. ""King of England"" he said ""The Red and White Knight on a Black and White Horse is here to see you"". The king turned to the guard and said ""Tell the Red and White Knight on a Black and White Horse that he may speak with me"".

The guard returned to the Red and White Knight on a Black and White Horse and said ""Red and White Knight on a Black and White Horse, the king has allowed you to see him, follow me"". 

So the Red and White Knight on a Black and White Horse followed the guard to the throne room and went and stood befor the king.

""Red and White Knight on a Black and White Horse what is it that you want from me"" said the King. The Red and White Knight on a Black and White Horse bowed before the king and said ""I the Red and White Knight on a Black and White Horse have come to ask for you daughters hand in Marriage"".

The king sat quietly to ponder the knights request for a few minutes and then said ""Red and White Knight on a Black and White Horse I will grant you my daughters hand in marriage if you get me the Shield of Glory from my Enemy the King of Wales"".

The red and white knight on a black and white horse replied ""I the Red and White Knight on a Black and White Horse will fetch you the sheild of Glory and then return for you daughter"".

The Red and White Knight on a Black and White Horse then left the castle and remounted on his trusty steed. 

The Red and White Knight on a Black and White Horse spent many weeks traveling to the King of Wales castle but finally arrived.

when he arrivd Red and White Knight on a Black and White Horse knocked on the gate of the king of Wales Castle. 

A few moments later a guard answered, he looked at the Red and White Knight on a Black and White Horse and said ""This is the castle of the king of wales who are you?"".

The Red and White Knight on a Black and White Horse got down off his horse and said ""I am the Red and White Knight on a Black and White Horse, and I want to see the King"" 

The guard looked at him for a while and said ""Red and White Knight on a Black and White Horse, I will ask the king if he will grant you an audience"".

The guard went through the castle and to the kings throne room. ""King of Wales"" he said ""The Red and White Knight on a Black and White Horse is here to see you"". The king turned to the guard and said ""Tell the Red and White Knight on a Black and White Horse that he may speak with me"".

The guard returned to the Red and White Knight on a Black and White Horse and said ""Red and White Knight on a Black and White Horse, the king has allowed you to see him, follow me"". 

So the Red and White Knight on a Black and White Horse followed the guard to the throne room and went and stood before the king.

""Red and White Knight on a Black and White Horse what is it that you want from me"" said the King. The Red and White Knight on a Black and White Horse bowed before the king and said ""I the Red and White Knight on a Black and White Horse have come to ask for you for the Sheild of Glory"".

The king sat quietly to ponder the knights request for a few minutes and then said ""Red and White Knight on a Black and White Horse I give you the Sheild of Glory If you get me the sword of might from my enemy the King of"".

The red and white knight on a black and white horse replied ""I the Red and White Knight on a Black and White Horse will fetch you the Sword of Might In exchange for the Sheild of Glory"".

The Red and White Knight on a Black and White Horse then left the castle and remounted on his trusty steed. 

The Red and White Knight on a Black and White Horse spent many weeks traveling to the King of Scotlands castle but finally arrived.

when he finally arrived the Red and White Knight on a Black and White Horse knocked on the gate of the king of Scotlands Castle. 

A few moments later a guard answered, he looked at the Red and White Knight on a Black and White Horse and said ""This is the castle of the king of Scotland who are you?"".

The Red and White Knight on a Black and White Horse got down off his horse and said ""I am the Red and White Knight on a Black and White Horse, and I want to see the King"" 

The guard looked at him for a while and said ""Red and White Knight on a Black and White Horse, I will ask the king if he will grant you an audience"".

The guard went through the castle and to the kings throne room. ""King of Scotland"" he said ""The Red and White Knight on a Black and White Horse is here to see you"". The king turned to the guard and said ""Tell the Red and White Knight on a Black and White Horse that he may speak with me"".

The guard returned to the Red and White Knight on a Black and White Horse and said ""Red and White Knight on a Black and White Horse, the king has allowed you to see him, follow me"". 

So the Red and White Knight on a Black and White Horse followed the guard to the throne room and went and stood before the king.

""Red and White Knight on a Black and White Horse what is it that you want from me"" said the King. The Red and White Knight on a Black and White Horse bowed before the king and said ""I the Red and White Knight on a Black and White Horse have come to ask for the sword of might"".

The king sat quietly to ponder the knights request for a few minutes and then said ""Red and White Knight on a Black and White Horse I will give you the sword of might if you fetch me the helm of power from my enemy the king of Ireland"".

The red and white knight on a black and white horse replied ""I the Red and White Knight on a Black and White Horse will fetch you the helm of power in exchange for the sword of might"".

The Red and White Knight on a Black and White Horse then left the castle and remounted on his trusty steed. 

The Red and White Knight on a Black and White Horse spent many weeks traveling to the King of Irelands castle but finally arrived.

One day the Red and White Knight on a Black and White Horse knocked on the gate of the king of Irelands Castle. 

A few moments later a guard answered, he looked at the Red and White Knight on a Black and White Horse and said ""This is the castle of the king of Ireland who are you?"".

The Red and White Knight on a Black and White Horse got down off his horse and said ""I am the Red and White Knight on a Black and White Horse, and I want to see the King"" 

The guard looked at him for a while and said ""Red and White Knight on a Black and White Horse, I will ask the king if he will grant you an audience"".

The guard went through the castle and to the kings throne room. ""King of Ireland"" he said ""The Red and White Knight on a Black and White Horse is here to see you"". The king turned to the guard and said ""Tell the Red and White Knight on a Black and White Horse that he may speak with me"".

The guard returned to the Red and White Knight on a Black and White Horse and said ""Red and White Knight on a Black and White Horse, the king has allowed you to see him, follow me"". 

So the Red and White Knight on a Black and White Horse followed the guard to the throne room and went and stood befor the king.

""Red and White Knight on a Black and White Horse what is it that you want from me"" said the King. The Red and White Knight on a Black and White Horse bowed before the king and said ""I the Red and White Knight on a Black and White Horse have come to ask for the Helm of Power"".

The king sat quietly to ponder the knights request for a few minutes and then said ""Red and White Knight on a Black and White Horse I will will give you my helm but only if you slay the Black and Blue Dragon with Green and Pink wings"".

The red and white knight on a black and white horse replied ""I the Red and White Knight on a Black and White Horse will slay the Black and Blue dragon with the green and pink wings"".

The Red and White Knight on a Black and White Horse then left the castle and remounted on his trusty steed. 

The Red and White Knight on a Black and White Horse travelled south to the lair of the Black and blue Dragon with the Green and pink wings.

After fighting for several days with the Black and Blue dragon with the Blue and Pink wings, The Red and White Knight on a Black and White horse finally slew the beast.

The Red and White Knight on a Black and White horse travelled all the way back to the King of Irelands castle.

When he arrived he knocked on the gate. A few minutes later the guard appeared. ""Red and White Knight on a Black and White horse, have you completed your quest?"".

The Red and White Knight on a Black and White horse replied ""I The Red and White Knight on a Black and White horse have defeated the Evil Black and Blue Dragon with the green and pink wings, and wish to see the king"".

""Follow me"" then said the guard, and he led The Red and White Knight on a Black and White horse to the kings throne room.

The king looked at The Red and White Knight on a Black and White horse and said ""Red and White Knight on a Black and White horse, have you slain the evil Black and blue Dragon with the Green and Pink wings?""

""Yes I The Red and White Knight on a Black and White horse have slain the dragon"" said the knight.

""Then here is the Helm of Power"" and the king gave the helm of power to The Red and White Knight on a Black and White horse.

The Red and White Knight on a Black and White horse left the Castle of the King of Ireland and and set off back to the king of scotlands Castle. 

When he arrived he knocked on the gate. A few minutes later the guard appeared. ""Red and White Knight on a Black and White horse, have you completed your quest?"".

The Red and White Knight on a Black and White horse replied ""I The Red and White Knight on a Black and White horse have the helm of power, and wish to see the king"".

""Follow me"" then said the guard, and he led The Red and White Knight on a Black and White horse to the kings throne room.

The king looked at The Red and White Knight on a Black and White horse and said ""Red and White Knight on a Black and White horse, have you got the helm of power?""

""Yes I The Red and White Knight on a Black and White horse have the helm of power.

""Then here is the sword of might"" and the king gave the sword of might to The Red and White Knight on a Black and White horse.

The Red and White Knight on a Black and White horse left the Castle of the King of scotland and and set off back to the king of wales Castle. 

When he arrived he knocked on the gate. A few minutes later the guard appeared. ""Red and White Knight on a Black and White horse, have you completed your quest?"".

The Red and White Knight on a Black and White horse replied ""I The Red and White Knight on a Black and White horse have the Sword of Might, and wish to see the king"".

""Follow me"" then said the guard, and he led The Red and White Knight on a Black and White horse to the kings throne room.

The king looked at The Red and White Knight on a Black and White horse and said ""Red and White Knight on a Black and White horse, do you have the Sword of might?""

""Yes I The Red and White Knight on a Black and White horse have the Sword of might.

""Then here is the Sheild of Glory"" and the king gave the Sheild of glory to The Red and White Knight on a Black and White horse.

The Red and White Knight on a Black and White horse left the Castle of the King of Wales and and set off back to the king of Englands Castle. 

When he arrived he knocked on the gate. A few minutes later the guard appeared. ""Red and White Knight on a Black and White horse, have you completed your quest?"".

The Red and White Knight on a Black and White horse replied ""I The Red and White Knight on a Black and White horse have the Sheild of Glory, and wish to see the king"".

""Follow me"" then said the guard, and he led The Red and White Knight on a Black and White horse to the kings throne room.

The king looked at The Red and White Knight on a Black and White horse and said ""Red and White Knight on a Black and White horse, Do you have the shield of Glory?""

""Yes I The Red and White Knight on a Black and White horse have slain the evil dragon to get the Helm of Power to get the Sword of Might to get the Shield of Glory, so can I now marry you daughter"".

And the King replied ""No"".",One day the Red and White Knight on a Black and White Horse knocked on the gate of the king of England's Castle.,0
post,4pudnd,2qh72,jokes,false,1466888537,https://old.reddit.com/r/Jokes/comments/4pudnd/im_naming_my_new_exercise_regime_brexit/,self.jokes,,It's the quickest way to lose pounds.,I'm naming my new exercise regime 'Brexit'.,11
post,4pudis,2qh72,jokes,false,1466888490,https://old.reddit.com/r/Jokes/comments/4pudis/a_hamburger_walks_into_a_bar/,self.jokes,,"Bartender says ""hey! We don't serve food here!""",A hamburger walks into a bar,139
post,4pudcb,2qh72,jokes,false,1466888415,https://old.reddit.com/r/Jokes/comments/4pudcb/my_wife_said_to_me_if_you_won_the_lottery_would/,self.jokes,,"I said: ""Of course I would. I'd miss you, but I'd still love you","My wife said to me: ""If you won the lottery, would you still love me?",200
post,4pud9w,2qh72,jokes,false,1466888391,https://old.reddit.com/r/Jokes/comments/4pud9w/hitlers_clone_was_just_found_out/,self.jokes,,[deleted],Hitler's clone was just found out...,0
post,4pud2t,2qh72,jokes,false,1466888320,https://old.reddit.com/r/Jokes/comments/4pud2t/how_many_lives_does_a_nazi_cat_have/,self.jokes,,"NEIN! 

I just realized that this actually makes sense because nein is the word for zero, and there aren't any Nazi cats (I mean they're all assholes, don't get me wrong, but they're not antisemitic). Multiple layers. Yay.",How many lives does a Nazi cat have?,1
post,4pucn6,2qh72,jokes,false,1466888167,https://old.reddit.com/r/Jokes/comments/4pucn6/aliens_finally_visit_earth/,self.jokes,,"Aliens suddenly show up on Earth.  They ask to meet with the world leaders, and as they greet each one, they hold up a small black rectangle up over their eyes for about 3 seconds and smile, then move on to greet the next.  After a while, one of the leaders asks, ""Why are you holding up the rectangle over your eyes?""

The aliens reply, ""We have been watching your species for several years, and whenever you come across another species from your planet, you do the same thing. We assumed it was the appropriate greeting."" The man is puzzled for a second but then remembers the smartphone in his pocket....",Aliens finally visit Earth...,0
post,4puciu,2qh72,jokes,false,1466888117,https://old.reddit.com/r/Jokes/comments/4puciu/a_poor_farmer_wants_a_vacation/,self.jokes,,"So he saves up money, then goes to a luxury hotel. The waiter gave him his key to his room, then told him where to go next. So the farmer did what he was told, but then a few minutes later, he stomped to the waiter, complaining:"" THAT IS A ROOM? YOU CAN'T EVEN PUT A CHAIR THERE! I'M OUT!"" 

The waiter laughed, then told the farmer: ""Sir, that's the elavator.""",A poor farmer wants a vacation.,6
post,4pucg1,2qh72,jokes,false,1466888091,https://old.reddit.com/r/Jokes/comments/4pucg1/a_man_goes_into_a_pharmacy/,self.jokes,,"A man goes into a pharmacy and buys a pack of condoms. As soon as he pays, he immediately starts laughing like a maniac and runs out of the pharmacy. The next day, the same man comes in, buys condoms, and runs out laughing. On the third day, when the man did it again, the pharmacist, a curious type by nature has his assistant follow the man. When the assistant comes back some time later, the pharmacists asks, ""so did you follow him?""

""Yes"" says the assistant

""And where did he go?"" 

""Home. Yours""",A man goes into a pharmacy,10
post,4puce9,2qh72,jokes,false,1466888072,https://old.reddit.com/r/Jokes/comments/4puce9/im_a_polish_student_in_the_uk/,self.jokes,,Today the cashier in ASDA asked me if I needed help packing my bags. The Brexit is worse than I thought...,I'm a Polish student in the UK,5
post,4pucbr,2qh72,jokes,false,1466888048,https://old.reddit.com/r/Jokes/comments/4pucbr/interviewer_where_do_you_see_yourself_in_10_years/,self.jokes,,[removed],Interviewer: where do you see yourself in 10 years? Me: in my clothes.,1
post,4pub9w,2qh72,jokes,false,1466887625,https://old.reddit.com/r/Jokes/comments/4pub9w/a_mans_car_breaks_down_in_a_blizzard_the_key_to/,self.jokes,,"John Jonson was making the yearly 400-mile-long trip to his relatives when snow began to fall. Small flakes, each intricate and delicate quickly turned to heavy gusts of snow. It didn't take long before John's vision was obscured and his car, to his dismay, began to cough and splutter. John, with his lack of mechanical knowledge, felt helplessly alone and scared. A man of 34, wife, kids, nice car, he never could have imagined he would die of anything other than old age, but the chill was creeping into his bones. A sudden feeling of determination to survive spurred John to pull down his cap, unbuckle his seat belt, and start a trek into the unknown to try to find shelter. Poor John lasted an admirable 20 minutes trekking before falling to his knees. Was this it? John thought. Will I never see my family again? 
     Just then, John saw a hand outstretched in front of him, offering help to his scrunched-up form. With closer inspection it was a man in simple orange garb, bare chest showing through his low V-necked robe. He wore no footwear, leading John to wonder how he could manage in the negative temperatures like that. The man lead him to a small, tucked away monastery in the hills. A roaring fire marked the end of a great hall; four hard wooden tables adorned with monks of all shapes and sizes. Simple wooden plates were filled with equally simple yet beckoning food, and John was happy to accept the offer of warmth and sustenance from the strange monks. 
      After a night of holy eating and conversing, John was led down a long hallway to his guest room. Sleeping for a few hours, he was suddenly awoken by the strangest sound. It's hard to put into words, like your classic, crackling, 'background noise' interspersed with sounds of birds and rushing water. John warily got out of bed and sheepishly opened his door, wandering down the long hall towards the sound. John's curiosity was rewarded when he came upon a huge, gold leaf adorned maple door, intricate and ornate, covered with strange letters the likes he had never seen before. The sound was much louder now; he felt strangely relaxed as it made its way in one ear and out of the other. After finding no door knob, John found his curiosity somewhat satiated, for now, and made his way back to a rewarding sleep. 
       In the morning, when John was eating breakfast with the 'head monk' who had helped him the night before, he asked him about the door. The monk replied 'I am sorry, young one, but I cannot tell you what is behind that door. You are not a monk.'. Gesturing to the tables of monks, he followed with 'We are welcoming to all, you may become a monk and see for yourself'. John hastily replied that he had a family, and did not mind too much.
       Happy to discover that the weather had cleared, and his car mysteriously fixed, John completed his trip, wondering about the strange door at first, but forgetting as he met with his family. 
       The next year, John was making the same trip, and at the *exact* same spot on the road as the last year, John broke down and a blizzard started whipping itself up. This time not hesitant, John stepped out of his car within a minute, and walked to where the monk had found him before. Lo and behold, the monk was standing in his spot. John made his way with his old friend to the tucked-away monastery, making friends with the new faces and once more going to bed, and slept. And again, he woke up after a few hours of disturbed sleep, to the other-worldly sound. Almost running down the corridor, he found himself before the mystical door, this time his entire body buzzing with spiritual energy. John made his way back to bed and slept once more.
In the morning, he asked the month just as he did last year, to *please* tell him what was behind the door. Rehearsed, the monk replied again 'I can't tell you, you're not a monk.'.
        Two years later, expecting it this time, John parked just before the blizzard and jogged to meet the monk. Excitedly, he told the monk that he was ready to become a monk! 'Very Good,' the monk said 'You shall know what you desire.'. 
           Ceremoniously, the monk led our protagonist down the long hall, knocking out a delicate yet deliberate beat against the door. Eager, John awaited a response. Nothing. Oh wait? What's this? The door, after seemingly eternity, finally started to creak open. Golden light shone out for a second, blinding John, and suddenly, as the light faded, he was exposed to what was beyond the door. Something so wondrous, people would kill to see it. Now, dear reader, would you like to see what John saw beyond the door?

 [I can't tell you, you're not a monk.](#s)",A man's car breaks down in a blizzard - the key to life,1
post,4pub5m,2qh72,jokes,false,1466887578,https://old.reddit.com/r/Jokes/comments/4pub5m/why_did_the_scarecrow_receive_an_award/,self.jokes,,[deleted],Why did the scarecrow receive an award?,0
post,4pu9ri,2qh72,jokes,false,1466887046,https://old.reddit.com/r/Jokes/comments/4pu9ri/you_matter/,self.jokes,,"Unless you multiply yourself by the speed of light squared.

Then you energy. ",You matter,6
post,4pu9i1,2qh72,jokes,false,1466886958,https://old.reddit.com/r/Jokes/comments/4pu9i1/how_do_you_stop_a_dog_from_humping_your_leg/,self.jokes,,... you pick him up and suck his dick.,How do you stop a dog from humping your leg?,4
post,4pu8za,2qh72,jokes,false,1466886767,https://old.reddit.com/r/Jokes/comments/4pu8za/what_do_the_amish_call_a_horse_with_gas/,self.jokes,,Air conditioning.,What do the Amish call a horse with gas?,1
post,4pu8p5,2qh72,jokes,false,1466886662,https://old.reddit.com/r/Jokes/comments/4pu8p5/son_i_want_you_to_give_this_letter_to_your_wife/,self.jokes,,[deleted],Son I want you to give this letter to your wife,0
post,4pu8ij,2qh72,jokes,false,1466886596,https://old.reddit.com/r/Jokes/comments/4pu8ij/hillary_clinton/,self.jokes,, ,Hillary Clinton,33
post,4pu8ay,2qh72,jokes,false,1466886512,https://old.reddit.com/r/Jokes/comments/4pu8ay/why_didnt_the_constipated_termite_become_a_doctor/,self.jokes,,[deleted],Why didn't the constipated termite become a doctor?,8
post,4pu7j4,2qh72,jokes,false,1466886186,https://old.reddit.com/r/Jokes/comments/4pu7j4/whos_got_the_biggest_list/,self.jokes,,Craig.,Who's got the biggest list?,0
post,4pu7ee,2qh72,jokes,false,1466886126,https://old.reddit.com/r/Jokes/comments/4pu7ee/why_cant_you_hear_a_pterodactyl_going_to_the/,self.jokes,,Because the P is silent.,Why can't you hear a pterodactyl going to the bathroom?,1
post,4pu70c,2qh72,jokes,false,1466885962,https://old.reddit.com/r/Jokes/comments/4pu70c/whats_the_hardest_part_about_eatting_a_vegetable/,self.jokes,,[deleted],What's the hardest part about eatting a vegetable?,2
post,4pu6vw,2qh72,jokes,false,1466885911,https://old.reddit.com/r/Jokes/comments/4pu6vw/hillary_clinton/,self.jokes,,[removed],Hillary Clinton.,1
post,4pu6k6,2qh72,jokes,false,1466885798,https://old.reddit.com/r/Jokes/comments/4pu6k6/johnnys_dad_said_do_your_revision/,self.jokes,,[deleted],"Johnny's dad said ""Do your revision!""",1
post,4pu6h2,2qh72,jokes,false,1466885764,https://old.reddit.com/r/Jokes/comments/4pu6h2/a_children_joking_with_teacher_amazing_you_can/,self.jokes,,[removed],A Children Joking With Teacher Amazing You Can Not Stop Laughing,1
post,4pu6ge,2qh72,jokes,false,1466885756,https://old.reddit.com/r/Jokes/comments/4pu6ge/whats_the_unforeseen_difference_ethernet_a_black/,self.jokes,,A snow tire doesn't sing when you put chai F sobe I t ,What's the unforeseen difference. Ethernet a black person and a snow tire.,0
post,4pu6ex,2qh72,jokes,false,1466885742,https://old.reddit.com/r/Jokes/comments/4pu6ex/a_family_is_at_the_dinner_table/,self.jokes,,"The father takes the chance to show off his new lie detecter robot that beeps when someone lies so he ask his son ""what we're you doing today son"" the son replies ""ummm I was at my friends house watching movies"" the robot beeps then the dad ask ""what we're you really doing son"" the son says guilty ""ok ok I was watching porn with my friend"" then the dad says ""I never watched porn when I was young"" the robot beeps and the mom says ""well that is your son"" the robot beeps",A family is at the dinner table,0
post,4pu65y,2qh72,jokes,false,1466885634,https://old.reddit.com/r/Jokes/comments/4pu65y/what_do_you_call_someone_who_photographs_fish/,self.jokes,,A school shooter,What do you call someone who photographs fish?,7
post,4pu5so,2qh72,jokes,false,1466885490,https://old.reddit.com/r/Jokes/comments/4pu5so/what_does_justin_timberlake_say_when_hes_going_to/,self.jokes,,"""It's Gonna Be Pee""",What does Justin Timberlake say when he's going to the bathroom?,0
post,4pu58y,2qh72,jokes,false,1466885263,https://old.reddit.com/r/Jokes/comments/4pu58y/how_can_jesus_prove_hes_holy/,self.jokes,,By holding up his hands. ,How can Jesus prove he's holy?,1
post,4pu4cg,2qh72,jokes,false,1466884918,https://old.reddit.com/r/Jokes/comments/4pu4cg/results_of_the_math_test_is_in/,self.jokes,,[deleted],Results of the math test is in,0
post,4pu485,2qh72,jokes,false,1466884868,https://old.reddit.com/r/Jokes/comments/4pu485/fun_presidential_trivia/,self.jokes,,"The annual salary of Commander-in-Chief is legally set at $400,000 per year. Except for our next one, who will only make $316,000 (or 79% to every man's dollar).",Fun Presidential Trivia,1
post,4pu37a,2qh72,jokes,false,1466884471,https://old.reddit.com/r/Jokes/comments/4pu37a/what_do_you_see_when_pillsbury_doughboy_bends_over/,self.jokes,,Donuts,What Do You See When Pillsbury Doughboy Bends Over?,19
post,4pu2kx,2qh72,jokes,false,1466884228,https://old.reddit.com/r/Jokes/comments/4pu2kx/britain_used_their_5050_and_ask_the_audience/,self.jokes,,"But it seems nobody understood it counts even if Chris Tarrant doesn't ask 'Is that your final answer?'

We should have used our bloody phone a friend.",Britain used their 50/50 and ask the audience.,0
post,4pu2k7,2qh72,jokes,false,1466884222,https://old.reddit.com/r/Jokes/comments/4pu2k7/id_tell_a_bondage_joke/,self.jokes,,But I'm all tied up.,I'd tell a bondage joke...,0
post,4pu2k6,2qh72,jokes,false,1466884222,https://old.reddit.com/r/Jokes/comments/4pu2k6/id_tell_a_bondage_joke/,self.jokes,,[deleted],I'd tell a bondage joke...,0
post,4pu2g0,2qh72,jokes,false,1466884182,https://old.reddit.com/r/Jokes/comments/4pu2g0/i_like_black_people_like_i_like_my_coffee/,self.jokes,,I don't like coffee.,I like black people like I like my coffee...,0
post,4pu1qw,2qh72,jokes,false,1466883901,https://old.reddit.com/r/Jokes/comments/4pu1qw/what_do_you_call_a_hip_arab/,self.jokes,,A chic sheik,What do you call a hip Arab?,0
post,4pu0wa,2qh72,jokes,false,1466883554,https://old.reddit.com/r/Jokes/comments/4pu0wa/a_train_owner_was_killed_by_a_wouldbe_engineer/,self.jokes,,Talk about a loco motive!,A train owner was killed by a would-be engineer over failing his operator's exam...,1
post,4pu0nm,2qh72,jokes,false,1466883463,https://old.reddit.com/r/Jokes/comments/4pu0nm/why_did_the_buddhist_businessman_have_more_money/,self.jokes,,[deleted],Why did the Buddhist businessman have more money?,0
post,4pu0fa,2qh72,jokes,false,1466883363,https://old.reddit.com/r/Jokes/comments/4pu0fa/i_have_a_joke/,self.jokes,,[deleted],I have a joke,0
post,4pu03a,2qh72,jokes,false,1466883234,https://old.reddit.com/r/Jokes/comments/4pu03a/i_told_my_gay_friend_i_could_turn_fruits_into/,self.jokes,,"He said ""prove it.""

So I pushed him off the balcony.",I told my gay friend I could turn fruits into vegetables...,1399
post,4ptzr2,2qh72,jokes,false,1466883104,https://old.reddit.com/r/Jokes/comments/4ptzr2/there_is_a_guy_who_always_wakes_up_surprised/,self.jokes,,One day he woke up and he wasn't surprised. So he got surprised!,There is a guy who always wakes up surprised.,1
post,4ptze7,2qh72,jokes,false,1466882971,https://old.reddit.com/r/Jokes/comments/4ptze7/i_get_pretty_nervous_when_my_phone_is_on_one_bar/,self.jokes,,It really puts me on Edge. ,I get pretty nervous when my phone is on one bar.,4
post,4ptz7f,2qh72,jokes,false,1466882902,https://old.reddit.com/r/Jokes/comments/4ptz7f/please_call_me_a_texi/,self.jokes,,[deleted],Please call me a texi,0
post,4ptyqs,2qh72,jokes,false,1466882731,https://old.reddit.com/r/Jokes/comments/4ptyqs/europe_classroom/,self.jokes,,"Classroom. All European Union countries are sitting. Britain raises a hand.  
-Teacher, Brussels, can I please leave?  
-Do you have a note from your nation? -the teacher inquires.  
-Yes, I do (Shows the note)  
-Oh, I see it has been written by your grandparents, well OK, you can go.

Someone is knocking the door, the doors open and there stands Ukraine asking to come in.  
Holland stands up saying ‘NO’.  
-Oh well - says Ukraine while closing the door - I will try later on.

Teacher Brussels says: 
-Ok, children, next week all of us are fundraising for the class to help sort the refugee crisis.   Germany rises a hand and says:  
-What? Is it again that everyone is meeting at mines? And why is it I have to pay the most for the fundraising.  
Brussell:  
-Here, everyone, look how well Germany is doing in the class. Always hands a helping hand, even when coming from a difficult family with a hard history… (looks at the back seats of the class) what about you there sitting at the back, Lithuania, Romania, Latvia… Are you going to take the example and become better students? How do you imagine your future?  
Lithuania from the back, while chewing on the sunflower seeds:  
- Eh.. It is fine, we can stay at someone’s from the class, like Ireland’s place.  
Ireland looks up:  
-Last time, you and Poland have stayed at mines, all of the silver was gone.

The door opens and Russia comes in.  
Brussels:  
-Oh, Russia, why did you not knock? Came in like it was your home.  
-Well, we are used to it (notices one empty seat). Oh, I see Britain have left the class. I will go tell my homeys, they will be happy",Europe Classroom,0
post,4pty99,2qh72,jokes,false,1466882544,https://old.reddit.com/r/Jokes/comments/4pty99/what_do_adolf_hitler_and_dale_earnhardt_have_in/,self.jokes,,[deleted],What do Adolf Hitler and Dale Earnhardt have in common?,0
post,4pty64,2qh72,jokes,false,1466882509,https://old.reddit.com/r/Jokes/comments/4pty64/so_the_president_of_nigeria_goes_to_russia/,self.jokes,,"When he arrives, he meets up with the president of Russia for a tour of the nation. ""I figured we could play a game that is *wildly* popular here, friend. It is called Russian roulette!""
The Nigerian president was curious, and asked how to play.
""Simple!"" said the Russian as he pulled out a revolver.
""you put *one bullet* into this gun, point it to your head, squeeze the trigger, and hope for the best.""
The Nigerian was no coward. He pulled the gun to his head after the Russian's succsesful attempt, and *click*
He was safe.
Weeks later, the Russian president paid a visit to his good friend in Nigeria.
He asked the Nigerian what their activities of the day would consist of. 
""My friend, today we play Nigerian roulette!""
The Nigerian clapped his hands and 6 beautiful women approached in front of the two men.
""Now here is how you play. Pick a woman, and she will give you the greatest blowjob you have *ever* had!""
The Russian was confused, and asked what the catch was.
The Nigerian laughed.
""You see my friend, one of these women happens to be a cannibal!""
",So the president of Nigeria goes to Russia..,117
post,4ptxvs,2qh72,jokes,false,1466882391,https://old.reddit.com/r/Jokes/comments/4ptxvs/why_did_the_chicken_cross_the_road/,self.jokes,,"TO GET TO THE OTHER SIDE!!!!


HahahahahahahahahahahahahahahahahahahahHAHAHAHAHAHAHAHAHAHAHAHAHHAHAHAHAHSHAHSHSGG OH....ohh...ha haha HAHAHAHHA HAHAHAHAHAHABHAA",wHy did the Chicken cross the road????,0
post,4ptxl3,2qh72,jokes,false,1466882280,https://old.reddit.com/r/Jokes/comments/4ptxl3/the_doctor_and_the_patient/,self.jokes,,"The doctor to the patient: 'You are very sick' 
The patient to the doctor: 'Can I get a second opinion?' 
The doctor again: 'Yes, you are very ugly too...'",The doctor and the patient,11
post,4ptx1o,2qh72,jokes,false,1466882072,https://old.reddit.com/r/Jokes/comments/4ptx1o/a_buddhist_monk_goes_to_a_barber/,self.jokes,,"..... to have his head shaved. ""What should I pay you?"" the monk asks. ""No price, for a holy man such as yourself,"" the barber replies. And what do you know, the next day the barber comes to open his shop, and finds on his doorstep a dozen gemstones.

That day, a priest comes in to have his hair cut. ""What shall I pay you, my son?"" ""No price, for a man of the cloth such as yourself."" And what do you know, the next day the barber comes to open his shop, and finds on his doorstep a dozen roses.

That day, Rabbi Finklestein comes in to get his payoss [sideburns] trimmed. ""What do you want I should pay you?"" ""Nothing, for a man of God such as yourself."" And the next morning, what do you know?

The barber finds on his doorstep — a dozen rabbis!
",A Buddhist monk goes to a barber,0
post,4ptwrf,2qh72,jokes,false,1466881961,https://old.reddit.com/r/Jokes/comments/4ptwrf/the_uk_is_dripping_more_pounds_than_jenny_craig/,self.jokes,,[removed],The UK is dripping more pounds than Jenny Craig,1
post,4ptwjv,2qh72,jokes,false,1466881875,https://old.reddit.com/r/Jokes/comments/4ptwjv/why_did_hitler_hate_the_jews/,self.jokes,,Because whenever he bought from them there was a high holocost,Why did Hitler hate the jews...,0
post,4ptvq5,2qh72,jokes,false,1466881562,https://old.reddit.com/r/Jokes/comments/4ptvq5/teacher_and_student/,self.jokes,,"Teacher: Whoever answers my next question, can go home. 

One boy throws his bag out the window. 

Teacher: Who just threw that? 

Boy: Me and I’m going home now.",Teacher and Student,305
post,4ptvgv,2qh72,jokes,false,1466881467,https://old.reddit.com/r/Jokes/comments/4ptvgv/aristotle_chipotle_i_rhyme_for_days_full_throttle/,self.jokes,,[deleted],"Aristotle, Chipotle, I rhyme for days full throttle",0
post,4ptvgs,2qh72,jokes,false,1466881465,https://old.reddit.com/r/Jokes/comments/4ptvgs/the_eyebrow_incident/,self.jokes,,[deleted],The Eyebrow Incident,1
post,4ptvg8,2qh72,jokes,false,1466881457,https://old.reddit.com/r/Jokes/comments/4ptvg8/breaking_news_oprah_arrested/,self.jokes,,"During a taping, police noticed something odd about her outfit. Upon searching, officers discovered 300 pounds of crack under her dress.",BREAKING NEWS: Oprah arrested!,0
post,4ptv4f,2qh72,jokes,false,1466881330,https://old.reddit.com/r/Jokes/comments/4ptv4f/a_man_decided_to_create_a_twitter_account_then/,self.jokes,,[deleted],A man decided to create a twitter account then deleted it...,0
post,4ptv3p,2qh72,jokes,false,1466881324,https://old.reddit.com/r/Jokes/comments/4ptv3p/doctor_patient_f/,self.jokes,,"Doctor: ""I'm sorry but you suffer from a terminal illness and have only 10 to live.""

Patient: ""What do you mean, 10? 10 what? Months? Weeks?!""

Doctor: ""Nine.""",Doctor &amp; Patient F,3
post,4ptuww,2qh72,jokes,false,1466881245,https://old.reddit.com/r/Jokes/comments/4ptuww/i_tried_suicide_once/,self.jokes,,I almost died :O,I tried suicide once,0
post,4ptust,2qh72,jokes,false,1466881197,https://old.reddit.com/r/Jokes/comments/4ptust/i_was_going_to_tell_a_joke_about_donald_trumps/,self.jokes,,"but then I realized it was racist,  too long, and didn't make any sense.",I was going to tell a joke about Donald Trump's presidential campaign..,8
post,4ptunk,2qh72,jokes,false,1466881136,https://old.reddit.com/r/Jokes/comments/4ptunk/at_school_we_were_always_taught_the_pullout/,self.jokes,,"...but like many teenagers, it hasn't stopped the UK trying anyway. ",At school we were always taught the pull-out method doesn't work...,144
post,4ptu95,2qh72,jokes,false,1466880967,https://old.reddit.com/r/Jokes/comments/4ptu95/im_surprised_that_the_uk_left_the_eu_by_voting/,self.jokes,,Most of the time they leave on penalty kicks.,I'm surprised that the UK left the EU by voting.,7
post,4ptu3l,2qh72,jokes,false,1466880906,https://old.reddit.com/r/Jokes/comments/4ptu3l/headline_leaves_eats_remains_for_brexit/,self.jokes,,[removed],Headline: Leaves Eats Remains for Brexit,1
post,4ptu1w,2qh72,jokes,false,1466880890,https://old.reddit.com/r/Jokes/comments/4ptu1w/im_a_call_you_chaps/,self.jokes,,Cause your sex life is assless.,I'm a call you Chaps...,0
post,4pttxt,2qh72,jokes,false,1466880840,https://old.reddit.com/r/Jokes/comments/4pttxt/what_happens_when_keemstar_and_ricegum_have_a_baby/,self.jokes,,He's born with Diss-lexia,What happens when Keemstar and Ricegum have a baby?,0
post,4pttn6,2qh72,jokes,false,1466880718,https://old.reddit.com/r/Jokes/comments/4pttn6/how_did_a_greet_b/,self.jokes,,[deleted],How did A greet B?,0
post,4pttft,2qh72,jokes,false,1466880644,https://old.reddit.com/r/Jokes/comments/4pttft/how_do_gay_people_make_coffee/,self.jokes,,[deleted],How do gay people make coffee?,0
post,4pttf3,2qh72,jokes,false,1466880635,https://old.reddit.com/r/Jokes/comments/4pttf3/i_cast_magic_missile_at_the_darkness/,self.jokes,https://www.reddit.com/r/Jokes/comments/4pttf3/i_cast_magic_missile_at_the_darkness/,,I cast magic missile at the darkness.,0
post,4ptsy5,2qh72,jokes,false,1466880449,https://old.reddit.com/r/Jokes/comments/4ptsy5/whats_the_difference_between_usain_bolt_and_adolf/,self.jokes,,Usain Bolt can finish a race.,What's the difference between Usain Bolt and Adolf Hitler?,69
post,4ptsnp,2qh72,jokes,false,1466880343,https://old.reddit.com/r/Jokes/comments/4ptsnp/since_yesterday_more_than_2_million_brits_have/,self.jokes,,That's what you get when Donald Trump says you made the right choice.,"Since yesterday, more than 2 million Brits have called for a new EU referendum...",6
post,4ptsgc,2qh72,jokes,false,1466880259,https://old.reddit.com/r/Jokes/comments/4ptsgc/what_does_a_sneeze_where_on_its_foot/,self.jokes,,[deleted],What does a sneeze where on its foot?,0
post,4pts5b,2qh72,jokes,false,1466880136,https://old.reddit.com/r/Jokes/comments/4pts5b/how_can_you_tell_if_a_person_is_a_vegetarian_in_a/,self.jokes,,"Don't worry, they WILL tell you.",How can you tell if a person is a vegetarian in a 5 minutes conversation?,0
post,4ptq5i,2qh72,jokes,false,1466879394,https://old.reddit.com/r/Jokes/comments/4ptq5i/what_do_you_call_a_country_that_leaves_the_eu/,self.jokes,,[deleted],What do you call a country that leaves the EU,0
post,4ptotc,2qh72,jokes,false,1466878876,https://old.reddit.com/r/Jokes/comments/4ptotc/nsfw_what_was_your_first_time_like/,self.jokes,,"Three friends are chilling in a bar, drinking and talking. One of them asks ""What was your first time like?"" 

The first guy says ""My first time was like riding a roller coaster. It started slow, then got really intense and fun, but it ended too quickly.""

The second guy says ""My first time was like watching a football game. I was having a blast, but she was so bored she was on her phone the entire time."" 

They both turn to look at the last guy, who sits quietly, thinking, until he finally speaks. ""My first time was like learning to ride a bicycle, with my dad holding my shoulders."" ","[NSFW] ""What was your first time like?""",42
post,4ptosz,2qh72,jokes,false,1466878874,https://old.reddit.com/r/Jokes/comments/4ptosz/mr_white_and_jesse_go_to_a_bar/,self.jokes,,[deleted],Mr White and Jesse go to a bar,0
post,4ptnnc,2qh72,jokes,false,1466878454,https://old.reddit.com/r/Jokes/comments/4ptnnc/whats_a_ghosts_favorite_type_of_music/,self.jokes,,Boograss!,What's a ghost's favorite type of music?,0
post,4ptn2c,2qh72,jokes,false,1466878243,https://old.reddit.com/r/Jokes/comments/4ptn2c/in_my_version_of_a_perfect_world_there_wouldnt_be/,self.jokes,,[deleted],"In my version of a perfect world, there wouldn't be any racism.",0
post,4ptmgv,2qh72,jokes,false,1466878019,https://old.reddit.com/r/Jokes/comments/4ptmgv/i_changed_my_bedding_as_a_gesture_of_hope/,self.jokes,,"I mean, if I can sheet the bed and have it work out, maybe the Brits can too.",I changed my bedding as a gesture of hope.,0
post,4ptmd5,2qh72,jokes,false,1466877974,https://old.reddit.com/r/Jokes/comments/4ptmd5/american_great/,self.jokes,,"I had to go see my doctor today because I’m having an unusual problem. I say to him, “I’ve got a problem, every time I finish masturbating I sing the American national anthem”.

The doctor said, “Don’t worry, a lot of wankers sing that”.",American great,6
post,4ptm5f,2qh72,jokes,false,1466877888,https://old.reddit.com/r/Jokes/comments/4ptm5f/did_you_hear_about_the_guy_who_didnt_accomplish/,self.jokes,,Neither did I.,Did you hear about the guy who didn't accomplish anything in his life?,3
post,4ptlar,2qh72,jokes,false,1466877572,https://old.reddit.com/r/Jokes/comments/4ptlar/why_is_it_hypocritical_of_the_republicans_to/,self.jokes,,[deleted],Why is it hypocritical of the Republicans to claim that creating a smaller government is their agenda?,0
post,4ptl5n,2qh72,jokes,false,1466877512,https://old.reddit.com/r/Jokes/comments/4ptl5n/3_men_are_stuck_on_an_island/,self.jokes,,"when they stumble upon a magic lamp. A genie comes out, and he says that he will give them each one wish. The first man says ""I wish to go home."" The second man says ""I wish to go home as well."" The third man says, ""I wish those other guys were back here, I'm lonely!""",3 men are stuck on an island...,0
post,4ptl0p,2qh72,jokes,false,1466877465,https://old.reddit.com/r/Jokes/comments/4ptl0p/a_man_heard_that_over_90_of_car_accidents_happen/,self.jokes,,So he moved.,A man heard that over 90% of car accidents happen within 15 km of home.,46
post,4ptk0y,2qh72,jokes,false,1466877059,https://old.reddit.com/r/Jokes/comments/4ptk0y/my_friend_said_he_knew_a_man/,self.jokes,,[removed],My friend said he knew a man,1
post,4ptjqp,2qh72,jokes,false,1466876945,https://old.reddit.com/r/Jokes/comments/4ptjqp/steam_summer_sale_2016_daily_deal_british_pound/,self.jokes,,[removed],Steam Summer sale 2016 daily deal! British Pound: 10% off,1
post,4ptjay,2qh72,jokes,false,1466876773,https://old.reddit.com/r/Jokes/comments/4ptjay/what_do_you_get_when_you_cross_stephen_colbert/,self.jokes,,John Oliver,What do you get when you cross Stephen Colbert with the entire country of England?,0
post,4ptjap,2qh72,jokes,false,1466876769,https://old.reddit.com/r/Jokes/comments/4ptjap/went_to_the_zoo_today/,self.jokes,,"I went to the zoo today, it sucked. Every thig was closed. They only had one animal. It was a shih tzu.",Went to the zoo today,0
post,4ptj7h,2qh72,jokes,false,1466876735,https://old.reddit.com/r/Jokes/comments/4ptj7h/why_do_cats_never_have_their_opinions_heard/,self.jokes,,"Because if it has a mu, it's not a statistic.",Why do cats never have their opinions heard?,1
post,4ptj3f,2qh72,jokes,false,1466876687,https://old.reddit.com/r/Jokes/comments/4ptj3f/whats_a_rappers_favorite_candy/,self.jokes,,Eminems.,What's a rapper's favorite candy?,4
post,4ptism,2qh72,jokes,false,1466876577,https://old.reddit.com/r/Jokes/comments/4ptism/what_do_we_call_rickon_stark/,self.jokes,,Plot device.,What do we call Rickon Stark?,0
post,4ptilk,2qh72,jokes,false,1466876498,https://old.reddit.com/r/Jokes/comments/4ptilk/the_eu/,self.jokes,,[deleted],The EU.,0
post,4ptij5,2qh72,jokes,false,1466876475,https://old.reddit.com/r/Jokes/comments/4ptij5/what_does_the_brazilian_pikachu_say/,self.jokes,,Zika zika.,What does the Brazilian Pikachu say?,72
post,4ptiew,2qh72,jokes,false,1466876427,https://old.reddit.com/r/Jokes/comments/4ptiew/jimmy_hendrix_eric_clapton_and_mick_jagger_are/,self.jokes,,"Jimmy trips over something in the sand and looks down to see a golden lamp. He picks it up and *POOF* out pops a genie. The genie looks at the men and says ""I will grant you each one wish for freeing me from the lamp!""

Hendrix goes first. ""I wish for a diamond the size of my head!"" He exclaims. The genie nods his head and *POOF* a huge diamond appears in Hendrix's hands.

Clapton gets excited and says, ""I wish for a massive yacht filled with beautiful women!"" The genie nods his head and *POOF* a yacht bigger than any they've ever seen pulls up to the Moroccan beach. 

The genie turns to Mick Jagger, who thinks for a minute, and finally says, ""I'm pretty hungry, I could go for a roll."" The genie nods his head and *POOF* a street vendor pushes his cart up the beach and hands Mick a delicious looking roll from his cart.

The genie vanishes and Hendix and Clapton give Jagger an incredulous look. ""You could have wished for anything in the world and that's what you wished for?!""

Jagger gives them a defensive look and says ""I know it's only a Moroccan roll, but I like it""  ","Jimmy Hendrix, Eric Clapton, and Mick Jagger are walking along the beach in Morocco...",15
post,4pthx6,2qh72,jokes,false,1466876239,https://old.reddit.com/r/Jokes/comments/4pthx6/what_do_you_call_a_cannibal_that_eats_relatives/,self.jokes,,Munchkin.,What do you call a cannibal that eats relatives?,11
post,4ptgfj,2qh72,jokes,false,1466875681,https://old.reddit.com/r/Jokes/comments/4ptgfj/last_time_i_was_this_early/,self.jokes,,[deleted],Last time I was this early...,0
post,4ptgcq,2qh72,jokes,false,1466875650,https://old.reddit.com/r/Jokes/comments/4ptgcq/an_elderly_couple_are_enjoying_their_75th/,self.jokes,,"The old man leans forward and says softly to his wife, “Dear, there is something that I must ask you. It has always bothered me that our tenth child never quite looked like the rest of our children. Now I want to assure you that these 75 years have been the most wonderful experience I could have ever hoped for, and your answer cannot take that all that away. But, I must know, did he have a different father?” The wife drops her head, unable to look her husband in the eye, she paused for a moment and then confessed. “Yes. Yes he did.” The old man is very shaken, the reality of what his wife was admitting hit him harder than he had expected. With a tear in his eye he asks “Who? Who was he? Who was the father?” Again the old woman drops her head, saying nothing at first as she tried to muster the courage to tell the truth to her husband. Then, finally, she says, “You.”",An elderly couple are enjoying their 75th anniversary.,453
post,4ptg2n,2qh72,jokes,false,1466875544,https://old.reddit.com/r/Jokes/comments/4ptg2n/why_do_trains_like_beef_jerky/,self.jokes,,[deleted],Why do trains like beef jerky?,0
post,4ptfun,2qh72,jokes,false,1466875461,https://old.reddit.com/r/Jokes/comments/4ptfun/whats_the_best_kind_of_cake_at_the_moment/,self.jokes,,Pound cake from the dollar store,What's the best kind of cake at the moment?,0
post,4ptet7,2qh72,jokes,false,1466875079,https://old.reddit.com/r/Jokes/comments/4ptet7/the_eu_now_has/,self.jokes,,[deleted],The EU now has..,0
post,4ptenj,2qh72,jokes,false,1466875013,https://old.reddit.com/r/Jokes/comments/4ptenj/a_guy_goes_to_the_supermarket_and_notices_an/,self.jokes,,[deleted],A guy goes to the supermarket and notices an attractive woman waving at him.,3
post,4ptdqu,2qh72,jokes,false,1466874664,https://old.reddit.com/r/Jokes/comments/4ptdqu/an_american_man_walks_into_a_bar/,self.jokes,,"An American man walks into a bar and as he sits down he overhears the conversation of the two women sitting next to him, speaking with British-sounding accents. He turns and asks, ""Excuse me ma'am, that's a lovely accent, are you women from England?"" The women instantly looked disgusted. One of them quickly and angrily replied ""Wales, you idiot!"" The man apologetically replied, ""I'm sorry, are you whales from England?""
",An American man walks into a bar...,1
post,4ptdd7,2qh72,jokes,false,1466874513,https://old.reddit.com/r/Jokes/comments/4ptdd7/my_mailman_got_gender_reassignment_surgery/,self.jokes,,Now he's a post man,My mailman got gender reassignment surgery.,520
post,4ptd5w,2qh72,jokes,false,1466874432,https://old.reddit.com/r/Jokes/comments/4ptd5w/oh_really/,self.jokes,,[removed],Oh really,0
post,4ptc3d,2qh72,jokes,false,1466874033,https://old.reddit.com/r/Jokes/comments/4ptc3d/whats_the_difference_between_adolf_hitler_and/,self.jokes,,Michael Schumacher can finish a race.,What's the difference between Adolf Hitler and Michael Schumacher?,1
post,4ptbz5,2qh72,jokes,false,1466873991,https://old.reddit.com/r/Jokes/comments/4ptbz5/limerick_there_once_was_a_man_from_waterloo/,self.jokes,,"A/N: This also works if you just say the first two lines out loud.
This joke may get you punched or called various names, for reasons soon apparent.

   
    There once was a man from Waterloo,
    whose limericks ended on line two.
        But that is such a bore,
        so this one ends line four.",[Limerick] There once was a man from Waterloo...,3
post,4ptbus,2qh72,jokes,false,1466873945,https://old.reddit.com/r/Jokes/comments/4ptbus/a_muslim_woman_came_to_the_husband_hajj/,self.jokes,,[deleted],A Muslim woman came to the husband Hajj,0
post,4ptbnd,2qh72,jokes,false,1466873861,https://old.reddit.com/r/Jokes/comments/4ptbnd/a_woman_goes_into_labour_and_her_husband_takes/,self.jokes,,"As she is laying in the hospital bed, the nurse tells her of a new type of technology that allows a percentage of her pain to be passed to the father of the child. They both agree, so start on 10% to be transferred.

However, the husband says he can feel nothing, and is willing for it to be turned up, so it goes up to 20%.

Again, he says the pain is bearable and more or less non-existent, so it goes up to 50%.

Eventually, the pain transfer gets turned up to 100%, and the husband is coping very well, allowing his wife to have a pain free child birth. ""This is so easy!"" he says.

Eventually, a healthy, adorable baby is born, and they get to take it home. They drive the whole way back smiling. They pull into their driveway and go to the front door, only to find the postman, dead on the doorstep.",A woman goes into labour and her husband takes her to the hospital.,995
post,4ptbgy,2qh72,jokes,false,1466873786,https://old.reddit.com/r/Jokes/comments/4ptbgy/dad_joke_lets_say_europe_has_caught_the_flu/,self.jokes,,[deleted],Dad joke: Let's say Europe has caught the flu...,1
post,4ptbfn,2qh72,jokes,false,1466873774,https://old.reddit.com/r/Jokes/comments/4ptbfn/the_turtle_lizard_and_rabbit/,self.jokes,,"One day, Turtle, Lizard, and Rabbit decide to start a garden. So as first things first they needed manure for their plants, Turtle and Lizard send the rabbit to town for the manure while they dig. While Rabbit was in town searching for the rich soil, Turtle and Lizard strike oil. As the rabbit returns he notices the rabbit and lizard are gone and there's a mansion where their farm was, so Rabbit knocks on the door and here comes a butler. Rabbit, confused as can be, asks the butler, where is Turtle and Lizard? The butler proceeds to say in a very classy tone, Mr. TurTEL is down by the well, and Mr. LizARD is near the yard. Then rabbit says, well you can tell them Mr.RabbIT is here with the shit!","The Turtle, Lizard, and Rabbit",1
post,4ptar6,2qh72,jokes,false,1466873487,https://old.reddit.com/r/Jokes/comments/4ptar6/the_us_drug_enforcement_agency_is_considering/,self.jokes,,Now there's a good iDEA,The US Drug Enforcement Agency is considering making an app for iPhone.,0
post,4pta9b,2qh72,jokes,false,1466873283,https://old.reddit.com/r/Jokes/comments/4pta9b/my_personal_favorite/,self.jokes,,[deleted],my personal favorite,3
post,4pta7e,2qh72,jokes,false,1466873262,https://old.reddit.com/r/Jokes/comments/4pta7e/why_was_the_tree_in_prison/,self.jokes,,because it committed treeson,Why was the tree in prison,18
post,4pt9ks,2qh72,jokes,false,1466873048,https://old.reddit.com/r/Jokes/comments/4pt9ks/an_englishman_a_scotsman_and_an_irishman_went_to/,self.jokes,,They all had to leave because the Englishman wanted to go.,"An Englishman, a Scotsman and an Irishman went to a bar.",1874
post,4pt9cd,2qh72,jokes,false,1466872962,https://old.reddit.com/r/Jokes/comments/4pt9cd/what_do_you_get_when_you_combine_two_japanese/,self.jokes,,A two-eyed onion.,What do you get when you combine two Japanese demons?,5
post,4pt8wo,2qh72,jokes,false,1466872805,https://old.reddit.com/r/Jokes/comments/4pt8wo/what_are_jewish_vampires_with_gluten_allergies/,self.jokes,,Garlic Nazis,What are Jewish vampires with gluten allergies most afraid of?,0
post,4pt8mz,2qh72,jokes,false,1466872701,https://old.reddit.com/r/Jokes/comments/4pt8mz/request_why_did_kamikaze_pilots_weared_helmets/,self.jokes,,[removed],[Request] Why did kamikaze pilots weared helmets?,1
post,4pt8bf,2qh72,jokes,false,1466872578,https://old.reddit.com/r/Jokes/comments/4pt8bf/2_whales/,self.jokes,,"2 whales walk into a bar.
First whale says: ooooEEEEEEEEaaaayyyyyuuuuuuaaaaaa eeeeooOOOOYAIIIAIIIEYOOOooooooo
Second whale says: Shut up Steve, you're drunk",2 whales,43
post,4pt832,2qh72,jokes,false,1466872490,https://old.reddit.com/r/Jokes/comments/4pt832/the_us_drug_enforcement_agency_is_considering/,self.jokes,,[deleted],The US Drug Enforcement Agency is considering making their own app,1
post,4pt82l,2qh72,jokes,false,1466872485,https://old.reddit.com/r/Jokes/comments/4pt82l/lance_armstrong/,self.jokes,,"I  think it is just terrible and disgusting how everyone has treated Lance Armstrong. Especially after what he achieved, winning 7 Tour de France races while on drugs. When I was on drugs, I couldn't even find my bike",Lance Armstrong,118
post,4pt7w3,2qh72,jokes,false,1466872419,https://old.reddit.com/r/Jokes/comments/4pt7w3/how_many_brits_does_it_take_to_change_a_broken/,self.jokes,,None. They just move out of the house.,How many Brits does it take to change a broken lightbulb?,526
post,4pt6vi,2qh72,jokes,false,1466872050,https://old.reddit.com/r/Jokes/comments/4pt6vi/what_do_you_call_the_area_where_a_horse_lives/,self.jokes,,The NEIGHHHHHHborhood,What do you call the area where a horse lives?,3
post,4pt6k7,2qh72,jokes,false,1466871935,https://old.reddit.com/r/Jokes/comments/4pt6k7/a_salesman_knocks_on_a_door/,self.jokes,,"It's answered by an eight-year-old wearing a smoking jacket. He has a scotch in one hand and a cigar in the other. 

Salesman says ""Hello young man, are your parents home?"". 

Kid says, ""Does it fucking look like it?"".",A salesman knocks on a door...,6
post,4pt68u,2qh72,jokes,false,1466871809,https://old.reddit.com/r/Jokes/comments/4pt68u/why_do_rogues_wear_leather_armoe/,self.jokes,,Because it's made of hide.,Why do rogues wear leather armoe?,45
post,4pt62l,2qh72,jokes,false,1466871734,https://old.reddit.com/r/Jokes/comments/4pt62l/this_referendum_is_getting_out_of_hand_now_wales/,self.jokes,,[removed],This Referendum Is getting out of hand. Now Wales and Northern Ireland are fighting!,1
post,4pt5id,2qh72,jokes,false,1466871514,https://old.reddit.com/r/Jokes/comments/4pt5id/small_dick_joke/,self.jokes,,Donald Trump,Small Dick Joke,0
post,4pt5c2,2qh72,jokes,false,1466871450,https://old.reddit.com/r/Jokes/comments/4pt5c2/a_man_walks_into_a_library_and_asks_for_a_book_on/,self.jokes,,[deleted],A man walks into a library and asks for a book on small penises,39
post,4pt4tq,2qh72,jokes,false,1466871260,https://old.reddit.com/r/Jokes/comments/4pt4tq/would_you_like_to_hear_a_story_about_my_friend/,self.jokes,,His name is Ali. Ali Gorical. ,Would you like to hear a story about my friend from Egypt?,0
post,4pt4e7,2qh72,jokes,false,1466871072,https://old.reddit.com/r/Jokes/comments/4pt4e7/i_dont_understand_why_people_think_donald_trump/,self.jokes,,[deleted],I don't understand why people think Donald Trump is making republicans look bad...,10
post,4pt49j,2qh72,jokes,false,1466871022,https://old.reddit.com/r/Jokes/comments/4pt49j/what_do_fall_out_boy_say_after_tittyfucking_their/,self.jokes,,THANKS FOR THE MAMMARIES!,What do Fall Out Boy say after titty-fucking their girlfriends?,3
post,4pt47t,2qh72,jokes,false,1466871006,https://old.reddit.com/r/Jokes/comments/4pt47t/like_my_uncle_used_to_say_the_best_part_of_twenty/,self.jokes,,...is there's twenty of them.,"Like my Uncle used to say, the best part of Twenty one year olds...",0
post,4pt468,2qh72,jokes,false,1466870989,https://old.reddit.com/r/Jokes/comments/4pt468/what_do_you_call_a_club_with_a_gun_range/,self.jokes,,[deleted],What do you call a club with a gun range?,0
post,4pt43x,2qh72,jokes,false,1466870964,https://old.reddit.com/r/Jokes/comments/4pt43x/whats_the_name_of_the_most_addicted_to_twitter/,self.jokes,,[deleted],What's the name of the most addicted to Twitter man in the world?,0
post,4pt3q6,2qh72,jokes,false,1466870808,https://old.reddit.com/r/Jokes/comments/4pt3q6/the_hairdressers/,self.jokes,,"Took my kid to the hairdressers the other day, she said ""aw your son has lovely curls"" I said ""yes he does"", She replied ""which side of the family does he get that from"", I said "" my friend has curly hair"".  ",The hairdressers,0
post,4pt32c,2qh72,jokes,false,1466870556,https://old.reddit.com/r/Jokes/comments/4pt32c/stalemate_on_four_letters/,self.jokes,,r/all,Stalemate on four (letters).,2
post,4pt2qy,2qh72,jokes,false,1466870430,https://old.reddit.com/r/Jokes/comments/4pt2qy/i_give_myself_an_excuse_for_watching_porn/,self.jokes,,"By pretending I'm watching ""How it's made: Babies"" on youtube.",I give myself an excuse for watching porn.,1
post,4pt25f,2qh72,jokes,false,1466870180,https://old.reddit.com/r/Jokes/comments/4pt25f/only_2000_kids_will_get_this/,self.jokes,,[deleted],Only 2000 kids will get this:,0
post,4pt25b,2qh72,jokes,false,1466870179,https://old.reddit.com/r/Jokes/comments/4pt25b/why_could_the_drunk_man_only_move_left/,self.jokes,,The officer hadn't read him his rights.,Why could the drunk man only move left?,9
post,4pt1ep,2qh72,jokes,false,1466869888,https://old.reddit.com/r/Jokes/comments/4pt1ep/how_do_you_keep_a_friend_in_suspense/,self.jokes,,[removed],How do you keep a friend in suspense?,1
post,4pt138,2qh72,jokes,false,1466869761,https://old.reddit.com/r/Jokes/comments/4pt138/the_uk_is_leaving_the_eu_and_because_of_that/,self.jokes,,So the english are going to get away scot free!,"The UK is leaving the EU and because of that, Scotland is moving for another Independence Referendum...",15
post,4pt0eu,2qh72,jokes,false,1466869496,https://old.reddit.com/r/Jokes/comments/4pt0eu/people_with_weight_problems/,self.jokes,,[deleted],People with weight problems...,8
post,4pt0ei,2qh72,jokes,false,1466869491,https://old.reddit.com/r/Jokes/comments/4pt0ei/hillary_clinton_is_elected_president/,self.jokes,,"On her first night in the White House (not counting when she was first lady), she is visited by the ghost of George Washington.

She asks, ""What can I do to help America?""

Washington replies ""Serve your country selflessly and always be honest""

*Hillary laughs in his face*

On her second day in the White House, she is visited by the ghost of Thomas Jefferson.

She asks, ""What can I do to help America?""

Jefferson replies ""Remember that governments derive their power from the consent of the governed, and that the individual is to have sovereignty over himself.""

*Hillary laughs in his face*

On her third day in the White House, she is visited by the ghost of Abraham Lincoln.

She asks, ""What can I do to help America?""

Lincoln replies ""Go to the theater.""",Hillary Clinton is elected President.,1171
post,4pt019,2qh72,jokes,false,1466869341,https://old.reddit.com/r/Jokes/comments/4pt019/a_man_was_going_hunting_with_his_friend/,self.jokes,,"While frantically tracking a wounded deer the men got separated.  In their haste to put the wounded animal out of its misery the man accidentally shot his friend in the chest, and his friend dropped with a thud.

Thankfully, he still had service in the woods and frantically dialed 911.  

""This is 911, what's your emergency?""

""I can't believe what happened!  I just shot my friend by accident while we were hunting, I think he's dead!""

""Ok sir please calm down. First make sure he's dead.""

The 911 operator waited for a moment and then a loud BANG was heard through the line.

""Okay, I'm sure he's dead.  Now what?""

",A man was going hunting with his friend.,15
post,4pszyu,2qh72,jokes,false,1466869309,https://old.reddit.com/r/Jokes/comments/4pszyu/how_many_twists_does_a_feminist_need_to_screw_in/,self.jokes,,None. They just grab it and the world to revolve around them.,How many twists does a feminist need to screw in a light bulb?,0
post,4pszae,2qh72,jokes,false,1466869036,https://old.reddit.com/r/Jokes/comments/4pszae/i_love_trump/,self.jokes,,[removed],I love Trump.,1
post,4psyvk,2qh72,jokes,false,1466868877,https://old.reddit.com/r/Jokes/comments/4psyvk/oh_that_seal/,self.jokes,,[removed],Oh that seal,1
post,4psysw,2qh72,jokes,false,1466868844,https://old.reddit.com/r/Jokes/comments/4psysw/what_did_god_say_to_mary_after_impregnating_her/,self.jokes,,Praise the Load,What did God say to Mary after impregnating her?,0
post,4psyro,2qh72,jokes,false,1466868833,https://old.reddit.com/r/Jokes/comments/4psyro/hey_theres_this_new_diet_that_can_help_lose/,self.jokes,,Its called the Brexit,Hey there's this new diet that can help lose pounds fast!,47
post,4psyqn,2qh72,jokes,false,1466868825,https://old.reddit.com/r/Jokes/comments/4psyqn/a_campfires_girlfriend_offers_to_give_him_a/,self.jokes,,[deleted],A campfire's girlfriend offers to give him a blowjob,0
post,4psykm,2qh72,jokes,false,1466868771,https://old.reddit.com/r/Jokes/comments/4psykm/teslas_are_so_safe_that_they_make_headlines_every/,self.jokes,,Probably because of the corduroy airbags,Teslas are so safe that they make headlines every time one crashes.,0
post,4psyjh,2qh72,jokes,false,1466868757,https://old.reddit.com/r/Jokes/comments/4psyjh/i_was_in_asda_and_then/,self.jokes,,"Just been to asda and there was a polish couple infront of me, the cashier said 'do you want help packing your bags?'                                       I thought bloody hell this is happening faster than i thought!",i was in asda and then...,0
post,4psxqo,2qh72,jokes,false,1466868448,https://old.reddit.com/r/Jokes/comments/4psxqo/the_eu_have_1_gb_free_space_now/,self.jokes,,[removed],The EU have 1 GB free space now,1
post,4psxik,2qh72,jokes,false,1466868344,https://old.reddit.com/r/Jokes/comments/4psxik/weird_computer_error/,self.jokes,,UK.eu has unexpectedly stopped working,Weird Computer Error,3
post,4pswye,2qh72,jokes,false,1466868092,https://old.reddit.com/r/Jokes/comments/4pswye/why_did_the_chicken_cross_the_road_nsfw/,self.jokes,,To suck the cock,Why did the chicken cross the road? (NSFW),0
post,4pswxg,2qh72,jokes,false,1466868084,https://old.reddit.com/r/Jokes/comments/4pswxg/i_lost_my_watch_at_a_party/,self.jokes,,"Saw a guy stepping on it while bullying a smaller dude. I walked up to the guy, and punched him. It's not okay to bully... not on my watch.",I lost my watch at a party...,85
post,4pswwb,2qh72,jokes,false,1466868076,https://old.reddit.com/r/Jokes/comments/4pswwb/brexit_slimming_product/,self.jokes,,"""Where can I get this new slimming product called ‪Brexit‬ ? I heard it helps you drop a lot of pounds.""",Brexit slimming product,0
post,4pswe0,2qh72,jokes,false,1466867869,https://old.reddit.com/r/Jokes/comments/4pswe0/i_guess_great_britain_is_going_for_its_roots/,self.jokes,,"Separated Kingdoms.
 

I'll see myself out.",I guess Great Britain is going for its roots...,1
post,4psw9z,2qh72,jokes,false,1466867823,https://old.reddit.com/r/Jokes/comments/4psw9z/now_that_britain_has_left_eu/,self.jokes,,Europe lost some storage space.. Exactly 1 GB ,Now that Britain has left EU,0
post,4psw41,2qh72,jokes,false,1466867762,https://old.reddit.com/r/Jokes/comments/4psw41/the_european_commission_has_just_announced_an/,self.jokes,,"As part of the negotiations, the British Government conceded that English spelling had some room for improvement and has accepted a 5- year phase-in plan that would become known as ""Euro-English"".


In the first year, ""s"" will replace the soft ""c"". Sertainly, this will make the sivil servants jump with joy. The hard ""c"" will be dropped in favour of ""k"". This should klear up konfusion, and keyboards kan have one less letter.

There will be growing publik enthusiasm in the sekond year when the troublesome ""ph"" will be replaced with ""f"". This will make words like fotograf 20% shorter.

In the 3rd year, publik akseptanse of the new spelling kan be expekted to reach the stage where more komplikated changes are possible.

Governments will enkourage the removal of double letters which have always ben a deterent to akurate speling.

Also, al wil agre that the horibl mes of the silent ""e"" in the languag is disgrasful and it should go away.

By the 4th yer people wil be reseptiv to steps such as replasing ""th"" with ""z"" and ""w"" with ""v"".

During ze fifz yer, ze unesesary ""o"" kan be dropd from vords kontaining ""ou"" and after ziz fifz yer, ve vil hav a reil sensi bl riten styl.

Zer vil be no mor trubl or difikultis and evrivun vil find it ezi TU understand ech oza. Ze drem of a united urop vil finali kum tru.
Und efter ze fifz yer, ve vil al be speking German like zey vunted in ze forst plas.

And Congratulations you have learnt German within minutes...","The European Commission has just announced an agreement whereby English will be the official language of the European Union rather than German, which was the other possibility.",22
post,4psv6h,2qh72,jokes,false,1466867383,https://old.reddit.com/r/Jokes/comments/4psv6h/what_tunnel_did_jews_go_through_the_most/,self.jokes,,The Chimney.,What tunnel did Jews go through the most?,0
post,4pstmw,2qh72,jokes,false,1466866746,https://old.reddit.com/r/Jokes/comments/4pstmw/the_english_language_will_now_only_have_3_vowels/,self.jokes,,"A, I, O.",The English language will now only have 3 vowels.,0
post,4pstiz,2qh72,jokes,false,1466866705,https://old.reddit.com/r/Jokes/comments/4pstiz/bad_roommate/,self.jokes,,"My college roommate from the past school year said that I was far better than his previous roommate. 
""He complained about me to the RA, and I constantly heard him fapping to porn,"" he recalled in disgust. ""When I used our bathroom after him, there would even be pubic hairs left on the edge of the sink.""
""What an asshole,"" I replied. ""I cleaned.""",Bad Roommate,0
post,4pstge,2qh72,jokes,false,1466866671,https://old.reddit.com/r/Jokes/comments/4pstge/eating_pistachios_is_like_picking_up_girls/,self.jokes,,You always go for the easiest ones to crack first.,Eating pistachios is like picking up girls,9
post,4pst2w,2qh72,jokes,false,1466866494,https://old.reddit.com/r/Jokes/comments/4pst2w/when_somebody_makes_you_really_angry_count_to/,self.jokes,,"When you get to two, punch them in the face. 

They won’t be expecting that.

","When somebody makes you really angry, count to three...",0
post,4pssyp,2qh72,jokes,false,1466866443,https://old.reddit.com/r/Jokes/comments/4pssyp/i_saw_a_girl_with_the_shortest_shorts_today/,self.jokes,,Her shorts were so short you could see private parts hanging out of mine!,I saw a girl with the shortest shorts today...,1
post,4pssy2,2qh72,jokes,false,1466866433,https://old.reddit.com/r/Jokes/comments/4pssy2/two_windmills_are_standing_in_a_field/,self.jokes,,"Two windmills are standing in a field and one asks the other, ""What kind of music do you like?""

The other says, ""I'm a big metal fan.""
",Two windmills are standing in a field...,0
post,4psskq,2qh72,jokes,false,1466866283,https://old.reddit.com/r/Jokes/comments/4psskq/ever_wonder_why_there_is_so_much_russian_anal_porn/,self.jokes,,[deleted],ever wonder why there is so much Russian anal porn?,1
post,4pssim,2qh72,jokes,false,1466866254,https://old.reddit.com/r/Jokes/comments/4pssim/i_put_a_dvd_on_ebay/,self.jokes,,6 people are watching it,I put a dvd on ebay,0
post,4pssbr,2qh72,jokes,false,1466866161,https://old.reddit.com/r/Jokes/comments/4pssbr/a_mans_wife_died_friend_asked_what_happend/,self.jokes,,"He said, she fell out from windows; as she was not drinking the poison. ",A man's wife died. friend asked what happend,0
post,4psrx7,2qh72,jokes,false,1466865978,https://old.reddit.com/r/Jokes/comments/4psrx7/what_do_you_call_a_dog_subbing_for_a_music_teacher/,self.jokes,,A subwoofer.,What do you call a dog subbing for a music teacher?,4
post,4psruw,2qh72,jokes,false,1466865953,https://old.reddit.com/r/Jokes/comments/4psruw/anti_joke_my_social_life/,self.jokes,,[deleted],Anti joke: my social life,5
post,4psru6,2qh72,jokes,false,1466865943,https://old.reddit.com/r/Jokes/comments/4psru6/i_read_a_joke_about_the_british_pound/,self.jokes,,But it didn't make any cents to me,I read a joke about the British pound...,5
post,4psqex,2qh72,jokes,false,1466865311,https://old.reddit.com/r/Jokes/comments/4psqex/the_united_states_and_britian_are_having_a/,self.jokes,,[deleted],The United States and Britian are having a competition on who can save Western Civilization.,0
post,4psqcn,2qh72,jokes,false,1466865283,https://old.reddit.com/r/Jokes/comments/4psqcn/two_immigrants_from_africa_arrive_in_the_united/,self.jokes,,"Two immigrants from Africa arrive in the United States and are discussing the difference between their country and the U.S. 

One of them mentions he's heard that people in the U.S. eat dogs, and if they're going to fit in, they better eat dogs as well. 

So they head to the nearest hot dog stand and order two 'dogs.' 

The first guy unwraps his, looks at it, and nervously looks at his friend. 

""Which part did you get?""

",Two immigrants from Africa arrive in the United States...,1429
post,4psp85,2qh72,jokes,false,1466864802,https://old.reddit.com/r/Jokes/comments/4psp85/how_many_brits_does_it_take_to_change_a_broken/,self.jokes,,[deleted],How many Brits does it take to change a broken lightbulb?,0
post,4psorv,2qh72,jokes,false,1466864575,https://old.reddit.com/r/Jokes/comments/4psorv/comedy_news_6_25_16/,self.jokes,,"Paul Ryan has an alternative to O'Bama-care. It involves the poor selling body parts &amp; a town crier yelling ""Bring out your dead""!

Hillary's slogan is 'I'm with her'. Wasn't that Chris Jenner's slogan as well?

I'll be performing at the world's largest music festival ""Summerfest"" on July 3rd at the Renegade Stage at 3 &amp; 5 :PM.

They're renovating the tomb of Jesus. How much upkeep foes that take? He was only there for 3 crummy days!

If I don't pay my bills, they turn off the electricity, cable, &amp; water. Doesn't that technically make me Amish? 

I'm on decaf now. That means I have no excuse for being a miserable jerk. I just have to learn to love myself even more.  

Good Humor has brought back it's ice cream trucks this summer. They're updated. They'll have armed guards &amp; sell ecstasy! 

My friend runs marathons for the 'runners high'. I'm so out of shape I get the same feeling if I stand up too quick!

They now have special 'kids menu's' at restaurants. Growing up the kids menu had 2 choices, 'eat it' or 'go hungry'! 


I'm planning my annual barbeque for July 9th. I like to schedule the first family fist fight between the potato salad and the baked beans. That leaves time to squeeze in the name calling &amp; threats before the watermelon!

",Comedy News 6 25 '16,1
post,4psop6,2qh72,jokes,false,1466864535,https://old.reddit.com/r/Jokes/comments/4psop6/the_united_states_and_britian_are_having_a/,self.jokes,,[deleted],The United States and Britian are having a competition on who can save the Western World.,0
post,4psob3,2qh72,jokes,false,1466864346,https://old.reddit.com/r/Jokes/comments/4psob3/how_did_tupac_die/,self.jokes,,[deleted],How did Tupac die?,0
post,4pso95,2qh72,jokes,false,1466864324,https://old.reddit.com/r/Jokes/comments/4pso95/why_did_the_chicken/,self.jokes,,[removed],Why did the chicken...,1
post,4pso34,2qh72,jokes,false,1466864242,https://old.reddit.com/r/Jokes/comments/4pso34/taking_a_shit/,self.jokes,,[deleted],Taking a Shit.,0
post,4pso1e,2qh72,jokes,false,1466864221,https://old.reddit.com/r/Jokes/comments/4pso1e/i_hope_england_beats_iceland/,self.jokes,,Or they will be out of Europe twice this week!,I hope England beats Iceland...,131
post,4psnnp,2qh72,jokes,false,1466864036,https://old.reddit.com/r/Jokes/comments/4psnnp/theres_that_moment_when_you_put_your_steak_on_the/,self.jokes,,"Do you vegans feel the same when you mow the grass?

",There’s that moment when you put your steak on the grill and your mouth waters all over from that amazing smell...,146
post,4psnj0,2qh72,jokes,false,1466863975,https://old.reddit.com/r/Jokes/comments/4psnj0/i_cant_wait_till_harriet_tubman_is_on_the_20_bill/,self.jokes,,That means I can legally own a black person again.,I can't wait till Harriet Tubman is on the $20 bill,0
post,4psmsd,2qh72,jokes,false,1466863618,https://old.reddit.com/r/Jokes/comments/4psmsd/there_are_three_unwritten_rules_of_life/,self.jokes,,[deleted],There are three unwritten rules of life:,1
post,4psl9r,2qh72,jokes,false,1466862873,https://old.reddit.com/r/Jokes/comments/4psl9r/why_do_girls_like_to_have_a_dog/,self.jokes,,"Because it suits their personality, a bitch.",Why do girls like to have a dog?,0
post,4psl5z,2qh72,jokes,false,1466862818,https://old.reddit.com/r/Jokes/comments/4psl5z/how_did_tupac_die/,self.jokes,,[deleted],How did Tupac die?,1
post,4psl30,2qh72,jokes,false,1466862780,https://old.reddit.com/r/Jokes/comments/4psl30/did_you_hear_about_the_guy_that_burned_off_his/,self.jokes,,The grease got so hot it caught fire when he tried to put it out it splashed up into his face burning his eyelids clean off. The doctors took his foreskin to make new eye lids. The procedure was a success but it left him a little cock-eyed.,Did you hear about the guy that burned off his eye lids in a kitchen fire?,1
post,4psk6i,2qh72,jokes,false,1466862333,https://old.reddit.com/r/Jokes/comments/4psk6i/this_one_might_be_a_little_over_the_top/,self.jokes,,[removed],This one might be a little over the top...,1
post,4psk3a,2qh72,jokes,false,1466862285,https://old.reddit.com/r/Jokes/comments/4psk3a/brexit_helped_me_with_my_weight_loss/,self.jokes,,I lost a bunch of pounds in a single day,Brexit helped me with my weight loss,0
post,4psjxu,2qh72,jokes,false,1466862210,https://old.reddit.com/r/Jokes/comments/4psjxu/taking_a_shit/,self.jokes,,[removed],Taking a shit,0
post,4psjv7,2qh72,jokes,false,1466862179,https://old.reddit.com/r/Jokes/comments/4psjv7/a_buddhist_monk_goes_to_a_barber_to_have_his_head/,self.jokes,," ""What should I pay you?"" the monk asks. ""No price, for a holy man such as yourself,"" the barber replies. And what do you know, the next day the barber comes to open his shop, and finds on his doorstep a dozen gemstones.


That day, a priest comes in to have his hair cut. ""What shall I pay you, my son?"" ""No price, for a man of the cloth such as yourself."" And what do you know, the next day the barber comes to open his shop, and finds on his doorstep a dozen roses.
 That day, Rabbi Finklestein comes in to get his payoss [sideburns] trimmed. ""What do you want I should pay you?"" ""Nothing, for a man of God such as yourself."" And the next morning, what do you know? The barber finds on his doorstep – a dozen rabbis
",A Buddhist monk goes to a barber to have his head shaved.,19918
post,4psiwt,2qh72,jokes,false,1466861668,https://old.reddit.com/r/Jokes/comments/4psiwt/today_brexit_helped_me_with_my_weight_loss/,self.jokes,,[deleted],Today Brexit helped me with my weight loss,1
post,4psiic,2qh72,jokes,false,1466861460,https://old.reddit.com/r/Jokes/comments/4psiic/whats_the_difference_between_donald_trump_and/,self.jokes,,[deleted],What's the difference between Donald Trump and Bitcoin?,0
post,4psi3f,2qh72,jokes,false,1466861261,https://old.reddit.com/r/Jokes/comments/4psi3f/i_tried_making_jokes_about_fat_people/,self.jokes,,... but none of them worked out.,I tried making jokes about fat people,60
post,4pshud,2qh72,jokes,false,1466861131,https://old.reddit.com/r/Jokes/comments/4pshud/what_does_a_siberian_kinkster_dream_of/,self.jokes,,[deleted],What does a Siberian kinkster dream of?,2
post,4psh90,2qh72,jokes,false,1466860817,https://old.reddit.com/r/Jokes/comments/4psh90/what_does_a_pirate_say_on_his_80th_birthday/,self.jokes,,[removed],What does a pirate say on his 80th birthday?,1
post,4psh30,2qh72,jokes,false,1466860738,https://old.reddit.com/r/Jokes/comments/4psh30/what_do_you_call_a_six_sided_shape_thats_missing/,self.jokes,,A hex-a-gone,What do you call a six sided shape that's missing?,30
post,4psgsm,2qh72,jokes,false,1466860591,https://old.reddit.com/r/Jokes/comments/4psgsm/its_no_wonder_germany_is_worried_about_brexit/,self.jokes,,"Last time they burned about a billion pounds, it didn't end well for them. ",It's no wonder Germany is worried about Brexit.,0
post,4psgez,2qh72,jokes,false,1466860404,https://old.reddit.com/r/Jokes/comments/4psgez/the_british_pound/,self.jokes,,[removed],The British Pound,1
post,4psfu4,2qh72,jokes,false,1466860135,https://old.reddit.com/r/Jokes/comments/4psfu4/i_have_just_finished_my_sandwich_degree/,self.jokes,, I do my final eggs ham tomorrow.,I have just finished my sandwich degree,1
post,4psf8i,2qh72,jokes,false,1466859830,https://old.reddit.com/r/Jokes/comments/4psf8i/i_got_fired_from_my_job_as_a_graphic_designer_my/,self.jokes,,[removed],I got fired from my job as a Graphic Designer. My work was too Graphic,1
post,4pseqy,2qh72,jokes,false,1466859575,https://old.reddit.com/r/Jokes/comments/4pseqy/disabled_toilets/,self.jokes,,"Ironically, the only toilets big enough to run around in.",Disabled toilets...,24
post,4psdzc,2qh72,jokes,false,1466859176,https://old.reddit.com/r/Jokes/comments/4psdzc/where_can_i_get_this_slimming_product_called/,self.jokes,,[deleted],Where can I get this slimming product called Brexit?,0
post,4psdt5,2qh72,jokes,false,1466859087,https://old.reddit.com/r/Jokes/comments/4psdt5/spoiler_what_is_hodors_favorite_band/,self.jokes,,The Doors.,[SPOILER] What is Hodor's favorite band?,0
post,4psdp1,2qh72,jokes,false,1466859025,https://old.reddit.com/r/Jokes/comments/4psdp1/the_european_union/,self.jokes,,[removed],The European Union,1
post,4psd3m,2qh72,jokes,false,1466858715,https://old.reddit.com/r/Jokes/comments/4psd3m/because_of_brexit/,self.jokes,,"James Bond is going to need a Visa for his Missions now. 
",Because of Brexit....,0
post,4pscjz,2qh72,jokes,false,1466858430,https://old.reddit.com/r/Jokes/comments/4pscjz/how_high_is_a_china_man_how_low_is_his_brother/,self.jokes,,[removed],How high is a China man How low is his brother,1
post,4psc72,2qh72,jokes,false,1466858271,https://old.reddit.com/r/Jokes/comments/4psc72/once_a_guy_needs_to_shit_very_badly/,self.jokes,,[deleted],once a guy needs to shit very badly,0
post,4psbrk,2qh72,jokes,false,1466858043,https://old.reddit.com/r/Jokes/comments/4psbrk/why_is_nobody_focusing_on_the_real_questions_of/,self.jokes,,like how are we going to tow the UK out of Europe?,Why is nobody focusing on the real questions of Brexit...,1
post,4psb5o,2qh72,jokes,false,1466857708,https://old.reddit.com/r/Jokes/comments/4psb5o/two_cows_walk_in_to_a_bar/,self.jokes,,"Then one of the cows says: ""*Mooooo*"", then the other replies,

""*Fuck, I was supposed to say that*""",Two cows walk in to a bar...,8
post,4psarj,2qh72,jokes,false,1466857467,https://old.reddit.com/r/Jokes/comments/4psarj/did_you_hear_about_the_incestuous_hotdogs/,self.jokes,,They say they're in bread. ,Did you hear about the incestuous hotdogs?,202
post,4psapv,2qh72,jokes,false,1466857438,https://old.reddit.com/r/Jokes/comments/4psapv/britain_leaving_the_eu_may_leave_a_rift_in_our/,self.jokes,,[deleted],Britain leaving the EU may leave a rift in our cultrues,0
post,4psakn,2qh72,jokes,false,1466857347,https://old.reddit.com/r/Jokes/comments/4psakn/give_me_some_gold/,self.jokes,,[deleted],Give me some gold...,0
post,4psag4,2qh72,jokes,false,1466857283,https://old.reddit.com/r/Jokes/comments/4psag4/a_dude_was_the_first_one_to_comment/,self.jokes,,"He said: ''Last time I was this early, the pound was still worth something''",A dude was the first one to comment.,2
post,4ps92r,2qh72,jokes,false,1466856492,https://old.reddit.com/r/Jokes/comments/4ps92r/nsfwbe_careful_what_you_wish_for/,self.jokes,,"A young man with a menial job was on his way home from work, and he finds an old lantern. Thinking that if he polishes it up he can get a few bucks for it.

He rubs the lamp and a genie comes out. The genie promises to grant him, three wishes.

Thinking he is on some reality TV show, he says Yeah right, but plays along.

He says to the genie, I wish I was rich, and the genie said granted. The man checks his bank balance and finds out that he is very rich.

Then the man says genie, I wish I was very handsome, and the genie said granted. The man pulls out a mirror and is astounded by how good he looks.

The man decides to save the wish for later, and the genie says that is fine, I will be listening.

The man goes home to decide what to do with his new found wealth and good looks.

He turns on the tv and there is an adult film playing. A buxom young woman is pleasuring herself with a large dildo. The man is turned on by the movie and says right now I wish I was a dildo, and the genie said granted.",[NSFW]Be careful what you wish for,0
post,4ps84y,2qh72,jokes,false,1466855985,https://old.reddit.com/r/Jokes/comments/4ps84y/for_women_life_is_a_lot_like_tetris/,self.jokes,,[deleted],"For women, life is a lot like tetris",23
post,4ps7q8,2qh72,jokes,false,1466855758,https://old.reddit.com/r/Jokes/comments/4ps7q8/whats_the_only_right_blacks_deserve/,self.jokes,,[removed],What's the only right blacks deserve?,0
post,4ps762,2qh72,jokes,false,1466855424,https://old.reddit.com/r/Jokes/comments/4ps762/good_news/,self.jokes,,[deleted],Good news!,0
post,4ps6g9,2qh72,jokes,false,1466855024,https://old.reddit.com/r/Jokes/comments/4ps6g9/how_come_arabs_are_not_circumcised/,self.jokes,,So they have some place to keep their gum safe during a sand storm. ,How come arabs are not circumcised?,0
post,4ps6fn,2qh72,jokes,false,1466855013,https://old.reddit.com/r/Jokes/comments/4ps6fn/trump/,self.jokes,,I wonder what would happen if Obama supported trump?,trump,0
post,4ps5zp,2qh72,jokes,false,1466854733,https://old.reddit.com/r/Jokes/comments/4ps5zp/so_i_was_walking_through_the_woods_and_i_came/,self.jokes,,[deleted],So i was walking through the woods and i came across a corpse,1
post,4ps5ul,2qh72,jokes,false,1466854642,https://old.reddit.com/r/Jokes/comments/4ps5ul/brexit_oxygen/,self.jokes,,[deleted],#Brexit &amp; oxygen,0
post,4ps5q5,2qh72,jokes,false,1466854556,https://old.reddit.com/r/Jokes/comments/4ps5q5/what_word_isnt_in_the_batdictionary/,self.jokes,,"Killing, unless your talking about his parents",What word isn't in the Bat-dictionary?,2
post,4ps5n5,2qh72,jokes,false,1466854493,https://old.reddit.com/r/Jokes/comments/4ps5n5/this_new_diet_is_great/,self.jokes,,[removed],This new diet is great!,1
post,4ps4nw,2qh72,jokes,false,1466853871,https://old.reddit.com/r/Jokes/comments/4ps4nw/the_only_reason_we_celebrate_our_birthdays/,self.jokes,,[deleted],The only reason we celebrate our birthdays,0
post,4ps4ks,2qh72,jokes,false,1466853817,https://old.reddit.com/r/Jokes/comments/4ps4ks/uk_votes_out_of_the_eu/,self.jokes,,[deleted],UK votes out of the EU...,0
post,4ps4ey,2qh72,jokes,false,1466853714,https://old.reddit.com/r/Jokes/comments/4ps4ey/last_time_i_got_some_ass/,self.jokes,,My finger went through the toilet paper,Last time I got some ass,10
post,4ps4at,2qh72,jokes,false,1466853625,https://old.reddit.com/r/Jokes/comments/4ps4at/have_you_seen_caitlyn_jenners_first_porno/,self.jokes,,[deleted],Have you seen Caitlyn Jenner's first porno?,0
post,4ps45w,2qh72,jokes,false,1466853527,https://old.reddit.com/r/Jokes/comments/4ps45w/whats_the_difference_between_a_dirty_bus_stop_and/,self.jokes,,"One's a crusty bus station, and one's a busty crustacean.",What's the difference between a dirty bus stop and a lobster with breast implants?,4
post,4ps44k,2qh72,jokes,false,1466853497,https://old.reddit.com/r/Jokes/comments/4ps44k/what_do_you_call_a_cow_with_no_legs/,self.jokes,,[deleted],What do you call a cow with no legs?,2
post,4ps3x0,2qh72,jokes,false,1466853369,https://old.reddit.com/r/Jokes/comments/4ps3x0/zoo/,self.jokes,,"I went to the zoo and saw a loaf in a cage.

A sign read: ""Bread in captivity.""",Zoo...,114
post,4ps3te,2qh72,jokes,false,1466853299,https://old.reddit.com/r/Jokes/comments/4ps3te/police_open_up/,self.jokes,," ""Police! Open up!""

 ""I don't want any balls!""

 ""We have no balls!""

 ""I know""","""Police! Open up!""",3
post,4ps3bu,2qh72,jokes,false,1466852994,https://old.reddit.com/r/Jokes/comments/4ps3bu/great_britains_new_prime_minister/,self.jokes,,Did you see that Boris Johnson might be the next Prime Minister of Great Britain? I remember when the U.S. had a BJ in the top office!,Great Britains new Prime Minister,13
post,4ps3bd,2qh72,jokes,false,1466852985,https://old.reddit.com/r/Jokes/comments/4ps3bd/what_do_you_call_a_person_eating_with_braces_on/,self.jokes,,[deleted],What do you call a person eating with braces on?,0
post,4ps35c,2qh72,jokes,false,1466852872,https://old.reddit.com/r/Jokes/comments/4ps35c/whats_an_arabs_favorite_car/,self.jokes,,Citroen C4,What's an Arab's favorite car?,0
post,4ps340,2qh72,jokes,false,1466852848,https://old.reddit.com/r/Jokes/comments/4ps340/uk_newspaper_headlines_yesterday_should_have_read/,self.jokes,,"EU referendum... EU sounds like 'you'. Thanks, I'll get my coat.

edit: changed al (Scots slang) to I'll... my bad Reddit, my bad!




","Uk newspaper headlines yesterday should have read as ""EU must be joking?!""",0
post,4ps2dd,2qh72,jokes,false,1466852365,https://old.reddit.com/r/Jokes/comments/4ps2dd/bob_told_his_wife_i_cant_work_for_him_anymore/,self.jokes,,"Wife: What did he say?

Bob: You're fired","Bob told his wife, ""I can't work for him anymore after what he said to me"".",329
post,4ps1vb,2qh72,jokes,false,1466852025,https://old.reddit.com/r/Jokes/comments/4ps1vb/my_grandfather_told_me_he_closed_one_eye_whenever/,self.jokes,,He was a sniper,My grandfather told me he closed one eye whenever he saw a jew in the good old days...,6
post,4ps1rq,2qh72,jokes,false,1466851953,https://old.reddit.com/r/Jokes/comments/4ps1rq/two_turds/,self.jokes,,[deleted],Two turds,1
post,4ps1ju,2qh72,jokes,false,1466851796,https://old.reddit.com/r/Jokes/comments/4ps1ju/tom_swifts_best_moments/,self.jokes,,"""German sausage jokes are the wurst,"" Tom said frankly.

""I got cut in half,"" Tom said intuitively.

""I will never read Shakespeare,"" Tom said unwillingly.

""I lost my legs right under the ankles,"" Tom said defeatedly.

""Who turned out the lights?"" Tom asked dimly.

""I don't know the words to this song,"" Tom said humbly.

""I lost my wrists,"" Tom said offhandedly.",Tom Swift's best moments.,10
post,4ps1by,2qh72,jokes,false,1466851653,https://old.reddit.com/r/Jokes/comments/4ps1by/as_you_can_see_the_eus_weight_loss_is_going_great/,self.jokes,,It lost all of its pounds.,As you can see the EU's weight loss is going great!,0
post,4ps0kx,2qh72,jokes,false,1466851167,https://old.reddit.com/r/Jokes/comments/4ps0kx/why_did_judy_hopps_find_it_difficult_to_rise_in/,self.jokes,,Because of the grass ceiling,Why did Judy Hopps find it difficult to rise in her career at the police department?,0
post,4ps0ap,2qh72,jokes,false,1466850991,https://old.reddit.com/r/Jokes/comments/4ps0ap/the_uk_must_be_taking_weight_loss_pills/,self.jokes,,[deleted],The UK must be taking weight loss pills...,2
post,4ps09m,2qh72,jokes,false,1466850971,https://old.reddit.com/r/Jokes/comments/4ps09m/my_dad_said_in_and_my_mum_said_out/,self.jokes,,[deleted],"My dad said ""in"" and my mum said ""out"".",0
post,4przo3,2qh72,jokes,false,1466850593,https://old.reddit.com/r/Jokes/comments/4przo3/all_these_brexit_jokes_are_getting_on_my_nerves/,self.jokes,,"I'm going to leave now.
",All these Brexit jokes are getting on my nerves..,0
post,4przf5,2qh72,jokes,false,1466850432,https://old.reddit.com/r/Jokes/comments/4przf5/mary_had_a_little_lamb/,self.jokes,,And also some orange juice to swallow it down with. ,Mary had a little lamb,0
post,4prz9m,2qh72,jokes,false,1466850328,https://old.reddit.com/r/Jokes/comments/4prz9m/someone_just_threw_a_bottle_of_omega_3_tablets_at/,self.jokes,,"I only suffered super fish oil injuries, but I'm lucky I wasn't krilled!




",Someone just threw a bottle of Omega 3 tablets at me.,32
post,4pryyq,2qh72,jokes,false,1466850144,https://old.reddit.com/r/Jokes/comments/4pryyq/what_happens_after_brexit/,self.jokes,,"Brexit could be followed by Grexit, Departugal, Italeave, Czechout, Oustria, Finish, Slovakout, Latervia and Byegium.  Looks like only Remania will stay..",What happens after Brexit.,0
post,4pryrp,2qh72,jokes,false,1466850013,https://old.reddit.com/r/Jokes/comments/4pryrp/latest_jobs_in_pakistan/,self.jokes,,[removed],Latest Jobs in Pakistan,1
post,4pryni,2qh72,jokes,false,1466849940,https://old.reddit.com/r/Jokes/comments/4pryni/i_like_putin/,self.jokes,,The rest of the joke down here,I like putin,49
post,4prw9b,2qh72,jokes,false,1466848390,https://old.reddit.com/r/Jokes/comments/4prw9b/whats_the_difference_between_a_black_man_and_a/,self.jokes,,The bench can support a family of four.,What's the difference between a black man and a bench?,1
post,4prvtw,2qh72,jokes,false,1466848120,https://old.reddit.com/r/Jokes/comments/4prvtw/i_think_britain_is_doing_quite_well_after_brexit/,self.jokes,,"In America, the bread bringer usually lose half his the assets after a divorce. Britain got off easy.",I think Britain is doing quite well after Brexit.,0
post,4prv0j,2qh72,jokes,false,1466847581,https://old.reddit.com/r/Jokes/comments/4prv0j/whats_the_difference_between_a_dirty_bus_stop_and/,self.jokes,,Ones a crusty bus station and ones a busty crustacean!,what's the difference between a dirty bus stop and a lobster with breast implants?,20
post,4pruk6,2qh72,jokes,false,1466847284,https://old.reddit.com/r/Jokes/comments/4pruk6/britain_can_now_say/,self.jokes,,...Its pull out game is strong!,Britain can now say....,9
post,4pruf5,2qh72,jokes,false,1466847184,https://old.reddit.com/r/Jokes/comments/4pruf5/this_brexit_thing_confuses_me/,self.jokes,,[deleted],This Brexit thing confuses me...,0
post,4pru8y,2qh72,jokes,false,1466847079,https://old.reddit.com/r/Jokes/comments/4pru8y/where_do_sex_offenders_go_after_death/,self.jokes,,[deleted],Where do sex offenders go after death?,3
post,4prtlu,2qh72,jokes,false,1466846609,https://old.reddit.com/r/Jokes/comments/4prtlu/if_minorities_have_the_race_card_women_have_the/,self.jokes,,[deleted],"If minorities have the race card, women have the gender card, and homosexuals have the gay card, what do discrimitory white men have?",1
post,4prspb,2qh72,jokes,false,1466845974,https://old.reddit.com/r/Jokes/comments/4prspb/the_captain_has_good_news_and_bad_news/,self.jokes,,"The Egyptian royal barge returns to harbour after a long day ferrying the pharaoh up and down the Nile. The captain says to the tired oarsmen 'Right, lads, I've got good news and bad news. Which do you want to hear first?'

The oarsmen consult among themselves and decide they fancy some good news first.

'The good news,' says the captain, 'Is that from now on your rations are doubled. The oarsmen cheer and start talking excitedly amongst themselves.

'The bad news,' says the captain, 'Is that Pharoah wants to try water-skiing.'",The captain has good news and bad news.,6
post,4prsi1,2qh72,jokes,false,1466845833,https://old.reddit.com/r/Jokes/comments/4prsi1/what_did_the_other_traffic_light_say_to_the_other/,self.jokes,,Don't look! I'm changing!,What did the other traffic light say to the other traffic light?,0
post,4prrw9,2qh72,jokes,false,1466845409,https://old.reddit.com/r/Jokes/comments/4prrw9/brexit_reform_bill_in_progress/,self.jokes,,[deleted],Brexit reform bill in progress...,3
post,4prr6e,2qh72,jokes,false,1466844902,https://old.reddit.com/r/Jokes/comments/4prr6e/i_wish_i_could_drop_pounds_as_fast_as_the_uk/,self.jokes,,[removed],I wish I could drop pounds as fast as the UK.,1
post,4prqzv,2qh72,jokes,false,1466844771,https://old.reddit.com/r/Jokes/comments/4prqzv/ive_recently_started_eating_steel/,self.jokes,,It's a refined taste,I've recently started eating steel,26
post,4prqoe,2qh72,jokes,false,1466844523,https://old.reddit.com/r/Jokes/comments/4prqoe/my_life/,self.jokes,,[removed],My life,1
post,4prqg6,2qh72,jokes,false,1466844348,https://old.reddit.com/r/Jokes/comments/4prqg6/i_was_in_tescos_yesterday/,self.jokes,,I was in tesco yesterday there was a Polish couple in front of me the lady at the check out asked if they needed help packing there bags I thought fucking hell love bit quick there,I was in tescos yesterday,6
post,4prpqh,2qh72,jokes,false,1466843854,https://old.reddit.com/r/Jokes/comments/4prpqh/man_sent_wife_to_buy_a_new_drill_gun/,self.jokes,,"... Worried for his wife, 2 hours later he gets a call from the police. ""Sir, you wife was arrested today, would you like to talk to her?"" Confused about what happened he said yes. ""What happened babe?!"" Wife says ""I just did what you asked, you told me to go to the store and find a black n decker""",Man sent wife to buy a new drill gun...,0
post,4prp3x,2qh72,jokes,false,1466843431,https://old.reddit.com/r/Jokes/comments/4prp3x/an_oldie_but_a_goodie/,self.jokes,,[removed],An oldie but a goodie!!,1
post,4prnu5,2qh72,jokes,false,1466842602,https://old.reddit.com/r/Jokes/comments/4prnu5/being_a_pornstar_must_be_the_best_job_ever/,self.jokes,,[deleted],Being a pornstar must be the best job ever...,0
post,4prnm6,2qh72,jokes,false,1466842470,https://old.reddit.com/r/Jokes/comments/4prnm6/how_high_is_a_china_man_how_low_is_his_brother/,self.jokes,,[removed],How high is a China man How low is his brother,1
post,4prnkl,2qh72,jokes,false,1466842441,https://old.reddit.com/r/Jokes/comments/4prnkl/a_black_family_ate_at_a_restaurant_and_tipped/,self.jokes,,[removed],A black family ate at a restaurant and tipped their server very well.,1
post,4prna0,2qh72,jokes,false,1466842230,https://old.reddit.com/r/Jokes/comments/4prna0/i_bought_a_llama_on_the_internet_today/,self.jokes,,[deleted],I bought a llama on the internet today.,1
post,4prn8n,2qh72,jokes,false,1466842207,https://old.reddit.com/r/Jokes/comments/4prn8n/its_easier_to_take_wales_out_of_the_eu/,self.jokes,,"...than it is to take a Welshman out of the ewe.
",It’s easier to take Wales out of the EU...,14
post,4prmkp,2qh72,jokes,false,1466841775,https://old.reddit.com/r/Jokes/comments/4prmkp/a_woman_walks_into_a_vet_with_her_duck/,self.jokes,,"It's being dragged behind her, evidently dead. She opens the door to an examining room and says ""I think my duck might be dead, doctor!"" The doctor says ""well ma'am, let me take a look"". So the doctor takes the duck and gently places it on the examining table. After a few quick checks, he says ""I'm sorry ma'am, your duck is dead"".

""That's impossible!"" She proclaims. ""I want a second opinion!"" So the doctor brings in a dog to confirm the finding. The dog sniffs the duck for a short while, then leaves the room. The doctor says ""I'm sorry ma'am, the dog concurs"". She is visibly upset now. She fights back tears and says ""are you absolutely sure, doctor?"" The doctor says ""well, we can check once more"".

So the doctor brings in a cat. The cat places its paws on the duck, pushes it a little, then walks out of the room, confirming that the duck is indeed dead. The woman, still clinging on to hope, says ""oh my, are you absolutely *certain*, doctor?"" The doctor replies ""yes ma'am, it was confirmed by myself, the lab results, and the cat scan"".",A woman walks into a vet with her duck,10
post,4prlyu,2qh72,jokes,false,1466841355,https://old.reddit.com/r/Jokes/comments/4prlyu/i_know_all_about_that/,self.jokes,,[removed],I know all about that...,0
post,4prl2o,2qh72,jokes,false,1466840759,https://old.reddit.com/r/Jokes/comments/4prl2o/what_do_you_get_when_you_cross_the_great_british/,self.jokes,,[deleted],What do you get when you cross the Great British Pound with BREXIT?,0
post,4prl0j,2qh72,jokes,false,1466840724,https://old.reddit.com/r/Jokes/comments/4prl0j/i_was_in_the_supermarket_today_and_the_cashier/,self.jokes,,"Fuck me, we only voted out yesterday give them a chance",I was in the supermarket today and the cashier asked the foreign couple in front of me if they needed help packing their bags,857
post,4prkm2,2qh72,jokes,false,1466840482,https://old.reddit.com/r/Jokes/comments/4prkm2/a_white_womans_waiting_in_line_at_the_grocery/,self.jokes,,[removed],A white woman's waiting in line at the grocery store...,0
post,4priq5,2qh72,jokes,false,1466839295,https://old.reddit.com/r/Jokes/comments/4priq5/little_johnny_once_bought_his_grandma_a_very_nice/,self.jokes,,"Little Johnny once bought his Grandma a very nice, luxurious toilet brush for her birthday. But when he went to visit her a couple of weeks later, it wasn't in the bathroom. 
Little Johnny asked his Grandma, “Gran, what happened to the toilet brush I gave you?”
“Darling, I'm sorry but I just didn’t like it. After all those years, I’ve gotten used to the toilet paper, and this new thing was just too scratchy.”",Little Johnny once bought his Grandma a very nice...,6
post,4pri8w,2qh72,jokes,false,1466838960,https://old.reddit.com/r/Jokes/comments/4pri8w/i_lost_my_mood_ring/,self.jokes,,I really just don't know how to feel about it. ,I lost my mood ring,19
post,4prfjx,2qh72,jokes,false,1466837333,https://old.reddit.com/r/Jokes/comments/4prfjx/the_pedophile_skipped_breakfast/,self.jokes,,[deleted],The pedophile skipped breakfast,0
post,4prf28,2qh72,jokes,false,1466837043,https://old.reddit.com/r/Jokes/comments/4prf28/when_i_eat_out_my_old_lady_you_know_what_she/,self.jokes,,[deleted],When I eat out my old lady you know what she tastes like?,0
post,4prezf,2qh72,jokes,false,1466836995,https://old.reddit.com/r/Jokes/comments/4prezf/the_british_currency_is_in_a_free_fall/,self.jokes,,"you can say it's gettin' pounded


[Please be gentle senpai.....it's my first time]",The British currency is in a free fall.....,0
post,4prele,2qh72,jokes,false,1466836772,https://old.reddit.com/r/Jokes/comments/4prele/whats_the_pounds_new_name/,self.jokes,,The ounce,What's the pound's new name?,3
post,4prdzx,2qh72,jokes,false,1466836434,https://old.reddit.com/r/Jokes/comments/4prdzx/a_little_boy_and_girl_are_talking/,self.jokes,,[deleted],A little boy and girl are talking...,5
post,4prdlw,2qh72,jokes,false,1466836209,https://old.reddit.com/r/Jokes/comments/4prdlw/a_string_walks_into_a_bar/,self.jokes,,"...and asks the bartender for a beer.
He nods toward a sign that says ""We don't serve strings!"". The string leaves and puts on a hat and walks back in. He tries to order a beer. The bartender goes to get one but looks at him suspiciously and asks ""Are you a string?"". The string says yes and leaves dejectedly. He makes one more effort and sneaks in through the bank door and goes into the bathroom. He ties the end of himself into a knot and frays the edges to look like hair. He goes to the bar and the bartender asks him....""Are you a string?""
The string replies....
""No, I'm a frayed knot!""",A string walks into a bar...,3
post,4prcc0,2qh72,jokes,false,1466835458,https://old.reddit.com/r/Jokes/comments/4prcc0/ever_wonder_why_britains_currency_dropped_so/,self.jokes,,Because paper money weighs like a gram but Britain's is a pound.,Ever wonder why Britain's currency dropped so quick after the Brexit compared to everyone else's?,2
post,4prbrt,2qh72,jokes,false,1466835144,https://old.reddit.com/r/Jokes/comments/4prbrt/genetic_link_to_obesity_proven/,self.jokes,,[removed],Genetic link to obesity proven,0
post,4prbor,2qh72,jokes,false,1466835096,https://old.reddit.com/r/Jokes/comments/4prbor/i_told_my_black_coworker_that_i_like_to_go_to/,self.jokes,,I said because I can't go to sleep listening to rap music and gunshots.,"I told my black coworker that I like to go to sleep listening to white noise. He said ""Why does it gotta be white noise with you people?""",42
post,4prbg8,2qh72,jokes,false,1466834963,https://old.reddit.com/r/Jokes/comments/4prbg8/the_rotation_of_the_earth/,self.jokes,,Really makes my day,The rotation of the earth,114
post,4prbg0,2qh72,jokes,false,1466834959,https://old.reddit.com/r/Jokes/comments/4prbg0/what_did_the_muslim_say_when_he_walked_into_the/,self.jokes,,[removed],What did the Muslim say when he walked into the bar?,0
post,4prb2i,2qh72,jokes,false,1466834737,https://old.reddit.com/r/Jokes/comments/4prb2i/what_do_you_call_a_school_with_majority_of_its/,self.jokes,,[removed],What do you call a school with majority of its students black?,0
post,4pram4,2qh72,jokes,false,1466834498,https://old.reddit.com/r/Jokes/comments/4pram4/i_was_going_to_use_the_new_machine_in_the_gym/,self.jokes,,But I found out it only sold protein bars,I was going to use the new machine in the gym,10
post,4pral6,2qh72,jokes,false,1466834487,https://old.reddit.com/r/Jokes/comments/4pral6/you_are_so_kind_funny_and_beautiful/,self.jokes,,"“Oh come on. You just want to get me to bed.” 


“And smart, too!","“You are so kind, funny and beautiful.”",1
post,4pra2f,2qh72,jokes,false,1466834219,https://old.reddit.com/r/Jokes/comments/4pra2f/a_muslim_man_walks_into_a_bar_and_says/,self.jokes,,[removed],A Muslim man walks into a bar and says...,1
post,4pr9a0,2qh72,jokes,false,1466833756,https://old.reddit.com/r/Jokes/comments/4pr9a0/how_can_you_make_number_seven_to_an_even_number/,self.jokes,,[deleted],How can you make number seven to an even number?,0
post,4pr8uq,2qh72,jokes,false,1466833522,https://old.reddit.com/r/Jokes/comments/4pr8uq/what_do_you_call_a_homosexual_on_roller_skates/,self.jokes,,[deleted],What do you call a homosexual on roller skates?,0
post,4pr8d7,2qh72,jokes,false,1466833281,https://old.reddit.com/r/Jokes/comments/4pr8d7/boss_hangs_a_poster_in_office/,self.jokes,,"Boss hangs a poster in office
‘I am the boss, dont forget’

He returns from lunch,
finds a slip on his desk,
‘ur wife called, she wants her poster back home..!!’",Boss hangs a poster in office,32
post,4pr8ca,2qh72,jokes,false,1466833270,https://old.reddit.com/r/Jokes/comments/4pr8ca/how_to_drink_a_coffee/,self.jokes,,"A customer ordered a cup of coffee in a restaurant! The waiter served the coffee. The customer found a fly in the coffee. He called the waiter.

Customer: How do I drink this coffee!
Waiter: Don’t you know how to drink a coffee? 
Customer: Waiter, see, there is a fly in my coffee. 
Waiter: Oh yes sir, you are right! There is a fly in your coffee. 
Customer: Waiter, I said, there is a fly in MMY coffee (He stressed the word MY)
Waiter: Oh don’t worry sir, the fly won’t drink much! 
Customer: Waiter, it is swimming in my coffee. 
Waiter: Sir, do you want me to get a lifeguard for the fly sir? 
(Annoyed) Customer: the fly dead, it’s irritating! 
Waiter: I guess, it doesn’t know how to swim properly. 
Customer: How do I drink this coffee? 
Waiter: Don’t you know how to drink? I will teach you! ",How to drink a coffee?,0
post,4pr840,2qh72,jokes,false,1466833145,https://old.reddit.com/r/Jokes/comments/4pr840/whats_the_opposite_of_a_gay_bar/,self.jokes,,An allahu akbar. ,What's the opposite of a gay bar?,1
post,4pr7h3,2qh72,jokes,false,1466832805,https://old.reddit.com/r/Jokes/comments/4pr7h3/longthe_turtle_lizard_and_rabbit/,self.jokes,,[deleted],"[Long]The Turtle, Lizard, and Rabbit",0
post,4pr79w,2qh72,jokes,false,1466832702,https://old.reddit.com/r/Jokes/comments/4pr79w/for_several_years_a_man_was_having_an_affair/,self.jokes,,"
with an Italian woman. One night, she confided in him that she was pregnant.
Not wanting to ruin his reputation or his marriage, he paid her a large sum of money if she would go to Italy to secretly have the child.
If she stayed in Italy to raise the child, he would also provide child support until the child turned 18. She tearfully agreed, but asked how to let him know when the baby was born.
To keep it discreet, he told her to simply mail him a postcard, and write “Spaghetti” on the back. He would then arrange for the child support payments to begin.
One day, about nine months later, he came home to his confused wife. “Honey,” she said, “you received a very strange postcard today.”
“Oh, just give it to me and I’ll explain it later,” he said.
The wife watched as her husband read the card, turned white, and fainted.

On the card was written:
“Spaghetti, Spaghetti, Spaghetti, Spaghetti, Spaghetti.
""Three with meatballs, two without. Send extra sauce.” ","For several years, a man was having an affair",202
post,4pr76f,2qh72,jokes,false,1466832656,https://old.reddit.com/r/Jokes/comments/4pr76f/just_overheard_the_funnest_conversation/,self.jokes,,[deleted],Just overheard the funnest conversation.,0
post,4pr6ty,2qh72,jokes,false,1466832478,https://old.reddit.com/r/Jokes/comments/4pr6ty/what_do_you_call/,self.jokes,,"what do you call a bunch of white people running down a hill?
-
-
-avalanche
what do you call a bunch of black people running down a hill?
-
-
-mudslide
what do you call a bunch of Mexicans running down a hill?
-
-
-jailbreak",what do you call.....,0
post,4pr6ki,2qh72,jokes,false,1466832347,https://old.reddit.com/r/Jokes/comments/4pr6ki/a_simple_way_to_lose_pounds_in_under_24_hours/,self.jokes,,Cut off your legs,A simple way to lose pounds in under 24 hours,8
post,4pr68k,2qh72,jokes,false,1466832160,https://old.reddit.com/r/Jokes/comments/4pr68k/cartunist/,self.jokes,,[deleted],Cartunist,0
post,4pr62j,2qh72,jokes,false,1466832061,https://old.reddit.com/r/Jokes/comments/4pr62j/two_nuns_are_driving_through_the_countryside_when/,self.jokes,,"The nun driving says to the passenger, ""Roll down the window and show him your cross!""

The other nun rolls down the window, leans out and shouts ""GET THE FUCK OFF OUR CAR!""","Two nuns are driving through the countryside, when a vampire jumps onto the roof of their car.",35
post,4pr61y,2qh72,jokes,false,1466832053,https://old.reddit.com/r/Jokes/comments/4pr61y/i_have_no_control_over_my_pasting/,self.jokes,,[removed],I have no control over my pasting.,1
post,4pr5t5,2qh72,jokes,false,1466831920,https://old.reddit.com/r/Jokes/comments/4pr5t5/boy_failed_to_reach_school_because_of_sign_on_the/,self.jokes,,[deleted],Boy failed to reach school because of Sign on the road,0
post,4pr5c1,2qh72,jokes,false,1466831672,https://old.reddit.com/r/Jokes/comments/4pr5c1/i_have_a_class_in_school_where_we_read_stories/,self.jokes,,It's lit,I have a class in school where we read stories and write reports on them.,1
post,4pr4fq,2qh72,jokes,false,1466831228,https://old.reddit.com/r/Jokes/comments/4pr4fq/which_one_is_closer_sun_or_africa/,self.jokes,,[deleted],"Which one is closer, Sun or Africa?",0
post,4pr3ux,2qh72,jokes,false,1466830931,https://old.reddit.com/r/Jokes/comments/4pr3ux/rocket_ship/,self.jokes,,"Did you hear about the rocket ship that didn't go up to space?

It had projectile dysfunction",Rocket Ship,4
post,4pr3u2,2qh72,jokes,false,1466830921,https://old.reddit.com/r/Jokes/comments/4pr3u2/european_union_has_lost_some_space/,self.jokes,,[deleted],European Union has lost some space,0
post,4pr3tq,2qh72,jokes,false,1466830917,https://old.reddit.com/r/Jokes/comments/4pr3tq/my_friend_told_me_that_recycling_is_good_for_the/,self.jokes,,"Not on Reddit, apparently. I got downvoted a lot...
",My friend told me that recycling is good for the environment,1
post,4pr3s9,2qh72,jokes,false,1466830896,https://old.reddit.com/r/Jokes/comments/4pr3s9/what_did_gandhi_fight_for/,self.jokes,,"Nothing, he was against violence.",What did Gandhi fight for?,0
post,4pr2kq,2qh72,jokes,false,1466830240,https://old.reddit.com/r/Jokes/comments/4pr2kq/i_had_my_wife_on_all_fours_last_night/,self.jokes,,As she was telling me to get out from under the bed and fight like a man. ,I had my wife on all fours last night...,25
post,4pr29q,2qh72,jokes,false,1466830060,https://old.reddit.com/r/Jokes/comments/4pr29q/a_polish_man_calls_911/,self.jokes,,"And says, ""Help! My wife is trying to kill me!""

The operator asks, ""How can you be sure?""

The Pole says, ""I was looking through her medicine cabinet, and I found Polish Remover!""",A Polish man calls 911,91
post,4pr1ez,2qh72,jokes,false,1466829604,https://old.reddit.com/r/Jokes/comments/4pr1ez/why_was_hitlers_suicide_such_a_suprise/,self.jokes,,Because we did nazi it coming,Why was hitler's suicide such a suprise?,0
post,4pr13m,2qh72,jokes,false,1466829457,https://old.reddit.com/r/Jokes/comments/4pr13m/theres_a_new_slimming_product_in_town_thatll_make/,self.jokes,,It's called brexit,There's a new slimming product in town that'll make you lose a lot of pounds,0
post,4pr0yo,2qh72,jokes,false,1466829388,https://old.reddit.com/r/Jokes/comments/4pr0yo/i_just_ate_a_frozen_apple/,self.jokes,,Hardcore.,I just ate a frozen apple!,11
post,4pr0ka,2qh72,jokes,false,1466829196,https://old.reddit.com/r/Jokes/comments/4pr0ka/why_did_the_pimps_garden_dry_up_and_die/,self.jokes,,Because all of his hose had kinks.,Why did the pimp's garden dry up and die?,0
post,4pr00c,2qh72,jokes,false,1466828913,https://old.reddit.com/r/Jokes/comments/4pr00c/why_is_india_surprised_by_the_brexit_vote/,self.jokes,,They didn't know you could get Britain to leave by voting.,Why is India surprised by the Brexit vote?,254
post,4pqzoz,2qh72,jokes,false,1466828752,https://old.reddit.com/r/Jokes/comments/4pqzoz/euna/,self.jokes,,[deleted],EU=NA?,0
post,4pqzex,2qh72,jokes,false,1466828607,https://old.reddit.com/r/Jokes/comments/4pqzex/finally_a_post_that_isnt_about_the_eu/,self.jokes,,So how about those Yankees?,Finally a post that isn't about the EU..,0
post,4pqxr8,2qh72,jokes,false,1466827786,https://old.reddit.com/r/Jokes/comments/4pqxr8/almost_got_raped_in_prison/,self.jokes,,My family takes Monopoly way too seriously,Almost got raped in prison,0
post,4pqxc0,2qh72,jokes,false,1466827578,https://old.reddit.com/r/Jokes/comments/4pqxc0/asking_for_a_pen/,self.jokes,,[deleted],Asking for a pen,0
post,4pqx65,2qh72,jokes,false,1466827505,https://old.reddit.com/r/Jokes/comments/4pqx65/mms/,self.jokes,,"Sometimes whenever I eat M&amp;Ms, I like to hold two M&amp;Ms in between my fingers and squeeze as hard as I can until one M&amp;M cracks, I eat the cracked one, and the one that didn't crack becomes the champion. Then I grab another M&amp;M and force it to compete with the champion in this deadly game of M&amp;M gladiators. I do this until I run out of M&amp;Ms and when there is only one M&amp;M left standing, I send a letter to M&amp;Ms brand with the champion M&amp;M in it with a note attached that reads: ""please use this M&amp;M for breeding purposes.""",M&amp;Ms,9
post,4pqx5z,2qh72,jokes,false,1466827502,https://old.reddit.com/r/Jokes/comments/4pqx5z/after_all_this_drama_with_the_brexit_maybe_if/,self.jokes,,[deleted],After all this drama with the Brexit. Maybe if Finland would leave ...,2
post,4pqwyy,2qh72,jokes,false,1466827411,https://old.reddit.com/r/Jokes/comments/4pqwyy/my_wife_punched_me_on_our_flight_from_georgia_to/,self.jokes,,[deleted],My wife punched me on our flight from Georgia to Kentucky.,0
post,4pqwx9,2qh72,jokes,false,1466827386,https://old.reddit.com/r/Jokes/comments/4pqwx9/why_is_moving_to_canada_always_plan_b/,self.jokes,,Canada deserves to be plan eh.,Why is moving to Canada always plan B?,2
post,4pqwbt,2qh72,jokes,false,1466827089,https://old.reddit.com/r/Jokes/comments/4pqwbt/a_man_was_having_a_horrible_day/,self.jokes,,[deleted],A man was having a horrible day...,9
post,4pqw2n,2qh72,jokes,false,1466826976,https://old.reddit.com/r/Jokes/comments/4pqw2n/if_gb_was_a_white_girl/,self.jokes,,European Union?!..... EU,If GB was a white girl...,0
post,4pqvb9,2qh72,jokes,false,1466826587,https://old.reddit.com/r/Jokes/comments/4pqvb9/a_man_is_walking_through_the_woods_when_he_comes/,self.jokes,,"Inside the suitcase he finds a fox and her cubs. He dials animal control to report his discovery. The woman on the other end exclaims, ""That's horrible... are they moving? The man responds, ""I don't know but that would explain the suitcase""",A man is walking through the woods when he comes across a suitcase.,1000
post,4pqv12,2qh72,jokes,false,1466826449,https://old.reddit.com/r/Jokes/comments/4pqv12/a_tree_tipped_over/,self.jokes,,A lot of pounds crashed to the ground,A tree tipped over,0
post,4pquse,2qh72,jokes,false,1466826329,https://old.reddit.com/r/Jokes/comments/4pquse/is_the_eu_working_out/,self.jokes,,It lost a few pounds this summer.,Is the EU working out?,7
post,4pqur1,2qh72,jokes,false,1466826309,https://old.reddit.com/r/Jokes/comments/4pqur1/whats_the_worst_thing_you_can_do_when_posting_a/,self.jokes,,Accidentally hit submit before you,What's the worst thing you can do when posting a joke?,7
post,4pqu7o,2qh72,jokes,false,1466826084,https://old.reddit.com/r/Jokes/comments/4pqu7o/did_you_hear_about_the_train_that_delivers_games/,self.jokes,,It's really picking up steam,Did you hear about the train that delivers games,11
post,4pqu2j,2qh72,jokes,false,1466826024,https://old.reddit.com/r/Jokes/comments/4pqu2j/the_united_states_and_britain_are_having_a/,self.jokes,,"Britain is in the lead, but America has a Trump card.",The United States and Britain are having a competition on who can fuck themselves up the most.,23359
post,4pqtmn,2qh72,jokes,false,1466825826,https://old.reddit.com/r/Jokes/comments/4pqtmn/what_is_nemos_favorite_kind_of_chip/,self.jokes,,Dory-tos           ;),What is Nemo's favorite kind of chip?,0
post,4pqsv1,2qh72,jokes,false,1466825471,https://old.reddit.com/r/Jokes/comments/4pqsv1/this_shark_was_teaching_his_kid_how_to_eat_humans/,self.jokes,,"He told him if you saw a human swimming,circle him 10 times and then attack

the kid looked to his father and said but why 10 times dad?

then the dad says well if you want to eat him with his shit go ahead",This shark was teaching his kid how to eat humans,5
post,4pqsr5,2qh72,jokes,false,1466825423,https://old.reddit.com/r/Jokes/comments/4pqsr5/my_friend_took_her_glasses_off/,self.jokes,,"The first thing my friend did is the cliche""how many fingers am I holding up?"" After she responded correctly, I asked her how many fingers God was holding up. She told me ""Allah dem""",My friend took her glasses off.,0
post,4pqre1,2qh72,jokes,false,1466824795,https://old.reddit.com/r/Jokes/comments/4pqre1/why_didnt_the_skeleton_cross_the_road/,self.jokes,,Why Didn't the skeleton cross the road? Because he didnt hav the guts :P,Why Didn't the skeleton cross the road?,3
post,4pqr5b,2qh72,jokes,false,1466824692,https://old.reddit.com/r/Jokes/comments/4pqr5b/any_love_for_trump_reversal_jokes/,self.jokes,,"In Obama's America, you serve the president, in Trump's America the president serves you. ",any love for Trump reversal jokes?,0
post,4pqr0j,2qh72,jokes,false,1466824628,https://old.reddit.com/r/Jokes/comments/4pqr0j/for_the_first_time_i_am_going_to_be_visiting/,self.jokes,,Britain had already left.,"For the first time I am going to be visiting Britain this summer, but when I got there...",3
post,4pqqs9,2qh72,jokes,false,1466824525,https://old.reddit.com/r/Jokes/comments/4pqqs9/one_day_scientists_will_make_a_very_powerful/,self.jokes,,[deleted],"One day, scientists will make a very powerful computer",2
post,4pqqp4,2qh72,jokes,false,1466824481,https://old.reddit.com/r/Jokes/comments/4pqqp4/what_is_et_shirt_for/,self.jokes,,It's because he has little legs ,What is ET shirt for?,0
post,4pqq9c,2qh72,jokes,false,1466824263,https://old.reddit.com/r/Jokes/comments/4pqq9c/how_do_you_cut_down_a_tree/,self.jokes,,A Suh dude,How do you cut down a tree?,0
post,4pqpzc,2qh72,jokes,false,1466824127,https://old.reddit.com/r/Jokes/comments/4pqpzc/what_did_the_lactose_intolerant_man_say_after/,self.jokes,,please excuse my dairy air ,what did the lactose intolerant man say after eating an ice cream cone?,6
post,4pqov1,2qh72,jokes,false,1466823626,https://old.reddit.com/r/Jokes/comments/4pqov1/donald_trump_has_written_a_lot_of_business_books/,self.jokes,,[deleted],Donald Trump has written a lot of business books.,4
post,4pqo4s,2qh72,jokes,false,1466823275,https://old.reddit.com/r/Jokes/comments/4pqo4s/why_was_hitler_so_robotic_and_nonsensical/,self.jokes,,[deleted],Why was Hitler so robotic and nonsensical?,0
post,4pqnlf,2qh72,jokes,false,1466823029,https://old.reddit.com/r/Jokes/comments/4pqnlf/i_have_sexdaily/,self.jokes,,I mean dyslexia fcuk,I have sexdaily,104
post,4pqnhv,2qh72,jokes,false,1466822984,https://old.reddit.com/r/Jokes/comments/4pqnhv/michael_jacksons_mom_was_recently_diagnosed_with/,self.jokes,,She had a bad mamma gramma,Michael Jackson's mom was recently diagnosed with Brest Cancer.,0
post,4pqngy,2qh72,jokes,false,1466822971,https://old.reddit.com/r/Jokes/comments/4pqngy/brexit_joke/,self.jokes,,The pound is rapidly losing value in currency exchange markets.,Brexit joke,0
post,4pqme3,2qh72,jokes,false,1466822522,https://old.reddit.com/r/Jokes/comments/4pqme3/why_were_hitlers_speeches_so_robotic_and/,self.jokes,,[deleted],Why were Hitler's speeches so robotic and nonsensical?,1
post,4pqlzk,2qh72,jokes,false,1466822335,https://old.reddit.com/r/Jokes/comments/4pqlzk/what_font_was_used_on_wyatt_earps_tombstone/,self.jokes,,Sans Sheriff.,What font was used on Wyatt Earp's tombstone?,15
post,4pqlre,2qh72,jokes,false,1466822240,https://old.reddit.com/r/Jokes/comments/4pqlre/i_dont_know_how_i_feel_about_masturbation_anymore/,self.jokes,,[deleted],I don't know how I feel about masturbation anymore...,7
post,4pqlqy,2qh72,jokes,false,1466822234,https://old.reddit.com/r/Jokes/comments/4pqlqy/why_do_all_of_the_drinks_in_vegas_and_hawaii_have/,self.jokes,,[deleted],why do all of the drinks in vegas and hawaii have straws?,0
post,4pqldh,2qh72,jokes,false,1466822080,https://old.reddit.com/r/Jokes/comments/4pqldh/what_did_the_tea_say_to_the_girl/,self.jokes,,[deleted],What did the tea say to the girl,0
post,4pqkpv,2qh72,jokes,false,1466821794,https://old.reddit.com/r/Jokes/comments/4pqkpv/if_donald_trump_becomes_president_and_boris/,self.jokes,,It'll be like toupees in a pod. ,"If Donald Trump becomes president, and Boris Johnson becomes UK's PM...",152
post,4pqkow,2qh72,jokes,false,1466821782,https://old.reddit.com/r/Jokes/comments/4pqkow/what_do_you_call_people_who_only_eat_vegetables/,self.jokes,,[deleted],What do you call people who only eat vegetables?,0
post,4pqkcs,2qh72,jokes,false,1466821643,https://old.reddit.com/r/Jokes/comments/4pqkcs/what_do_you_call_jokes_about_the_brexit/,self.jokes,,Branter.,What do you call jokes about the Brexit?,0
post,4pqkai,2qh72,jokes,false,1466821617,https://old.reddit.com/r/Jokes/comments/4pqkai/raw_egg_yokes_build_muscle/,self.jokes,,[deleted],Raw Egg Yokes Build Muscle,2
post,4pqkaa,2qh72,jokes,false,1466821614,https://old.reddit.com/r/Jokes/comments/4pqkaa/what_font_was_used_on_wyatt_earps_tombstone/,self.jokes,,[deleted],What font was used on Wyatt Earp's tombstone?,1
post,4pqjsr,2qh72,jokes,false,1466821375,https://old.reddit.com/r/Jokes/comments/4pqjsr/google_reports_consistent_level_of_searches_for/,self.jokes,,Title,"Google reports consistent level of searches for ""pornography"" in the UK following Brexit",0
post,4pqjdx,2qh72,jokes,false,1466821179,https://old.reddit.com/r/Jokes/comments/4pqjdx/in_the_old_days_folks_used_to_say_tisk_tisk_to/,self.jokes,,"Now social media connects us to millions, and allows us to multi-tisk. ","In the old days, folks used to say ""tisk, tisk"" to shame others",8
post,4pqj7a,2qh72,jokes,false,1466821100,https://old.reddit.com/r/Jokes/comments/4pqj7a/jews_be_like/,self.jokes,,[deleted],Jews be like...,0
post,4pqhyt,2qh72,jokes,false,1466820531,https://old.reddit.com/r/Jokes/comments/4pqhyt/the_secret_to_losing_pounds_in_less_than_24_hours/,self.jokes,,[deleted],The secret to losing pounds in less than 24 hours?,7
post,4pqhhb,2qh72,jokes,false,1466820324,https://old.reddit.com/r/Jokes/comments/4pqhhb/where_do_you_find_a_man_with_an_aquatic_mammal/,self.jokes,,In Wales.,Where do you find a man with an aquatic mammal fetish?,91
post,4pqhfj,2qh72,jokes,false,1466820302,https://old.reddit.com/r/Jokes/comments/4pqhfj/it_was_hard_until_i_came_into_faith_and_found/,self.jokes,,She was kind of pissed when she realized I wasn't using a condom though...,It was hard until I came into Faith and found bliss,4
post,4pqgwk,2qh72,jokes,false,1466820062,https://old.reddit.com/r/Jokes/comments/4pqgwk/the_stock_market_has_been_looking_thinner_lately/,self.jokes,,It's lost several Pounds.,The stock market has been looking thinner lately.,2
post,4pqgns,2qh72,jokes,false,1466819951,https://old.reddit.com/r/Jokes/comments/4pqgns/whats_the_difference_between_manual_driving_and/,self.jokes,,"Automatic driving is like having sex with a woman, It's natural and pretty enjoyable.

Manual driving is like having sex with a dude, a huge pain in the ass and you gotta handle the shaft most of the time, and disturbingly, some people begin to like it.

",What's the difference between manual driving and automatic driving?,0
post,4pqgls,2qh72,jokes,false,1466819929,https://old.reddit.com/r/Jokes/comments/4pqgls/what_does_a_scotsman_wear_under_his_kilt/,self.jokes,,Shame and sadness at the slow decline of their once beautiful and vibrant culture.,What does a Scotsman wear under his kilt?,2
post,4pqgka,2qh72,jokes,false,1466819910,https://old.reddit.com/r/Jokes/comments/4pqgka/a_chinese_family_moved_into_my_neighborhood_when/,self.jokes,,"They had a pair of twins, named Ving and Ling, who were my age. I liked Ving, but his sister Ling was kind of a bitch. Eventually, Ling told me that he hated his name, and he wanted to change it. I asked him, ""What do you want to change your name to?"" and he said ""Lee. You know, like Bruce Lee?"" Ling overheard, and chimed in, saying that their father would disown him if he changed his name.

One day, Ving decided he had had enough. He went to town hall, with me in tow. His sister caught wind and decided to come along  to talk him out of it. 

So we got the name change document, and Ving filled it out and almost turned it in, when he suddenly got choked up and realized that he couldn't go through with the name change. He told the receptionist that he wanted to cancel, and she told him that he could cancel the name change, but he'd need to pay a one-time fee of $20. Ving didn't have any money on him, but his sister did. She was about to hand him $20 when suddenly, a short, elderly Chinese man in an American flag T-shirt, ray-bans and cargo shorts entered the building. Ving stared at him in awe.

""D..Dad?"" he stammered, tearfully. 

With a huge smile on his face, the man ran up and embraced his son.

I'll never forget what his father said that day:

&gt; ""Don't stop, be Lee, Ving.  
&gt; Hold on the that fee, Ling""",A Chinese family moved into my neighborhood when I was in high school...,504
post,4pqg7x,2qh72,jokes,false,1466819751,https://old.reddit.com/r/Jokes/comments/4pqg7x/hey_girl_are_you_the_european_union/,self.jokes,,Because I don't know what you are or what you do but I am out of here. ,Hey Girl are you the European Union?,0
post,4pqfwv,2qh72,jokes,false,1466819606,https://old.reddit.com/r/Jokes/comments/4pqfwv/i_heard_brits_want_to_move_to_canada/,self.jokes,,[deleted],I heard Brits want to move to Canada,8
post,4pqfgy,2qh72,jokes,false,1466819423,https://old.reddit.com/r/Jokes/comments/4pqfgy/how_do_you_tell_if_a_man_is_gay/,self.jokes,,"When you're fucking him in the ass, reach around; if he has a boner... He's gay ",How do you tell if a man is gay?,27
post,4pqfc5,2qh72,jokes,false,1466819353,https://old.reddit.com/r/Jokes/comments/4pqfc5/what_do_you_call_a_gossiping_mushroom/,self.jokes,,[deleted],What do you call a gossiping mushroom?,14
post,4pqen5,2qh72,jokes,false,1466819049,https://old.reddit.com/r/Jokes/comments/4pqen5/what_did_the_doctor_say_to_the_obese_patient/,self.jokes,,It is time you lose a few pounds!,What did the doctor say to the obese patient after Brexit?,0
post,4pqe88,2qh72,jokes,false,1466818868,https://old.reddit.com/r/Jokes/comments/4pqe88/a_tale_of_two_photos/,self.jokes,,"A solider out at war, missing his mother and his girlfriend, decided to take a couple of pictures of himself to send to them. For his mother, he dressed up real nice and took a picture of himself from the torso up. For his girlfriend, he decided to take a picture of his nether regions. The solider then took the photos to the post office to be sent out. Unfortunately the photos got switched while sending, and so the girlfriend and the mother received the opposite photos.

When the girlfriend received the photo of her sharply-dressed man, she responded with ""Oh my, he looks so handsome!""

The mother, on the other hand, was old and fairly blind. Upon receiving the picture of her son, she became slightly upset. Taking a good look at the photo, she responded with ""Oh, my poor soon! It looks like he hasn't shaved in months! And his tie looks a bit crooked too...""",A Tale of Two Photos,8
post,4pqe1o,2qh72,jokes,false,1466818786,https://old.reddit.com/r/Jokes/comments/4pqe1o/coming_soon_to_the_usa/,self.jokes,, #Mexit,Coming soon to the USA...,3
post,4pqe0m,2qh72,jokes,false,1466818774,https://old.reddit.com/r/Jokes/comments/4pqe0m/if_orange_is_the_new_black/,self.jokes,,then Donald Trump is black,If orange is the new black?,2
post,4pqd8r,2qh72,jokes,false,1466818448,https://old.reddit.com/r/Jokes/comments/4pqd8r/silence_is_the_best_response_to_a_fool/,self.jokes,,[removed],Silence is the best response to a fool.,0
post,4pqcp0,2qh72,jokes,false,1466818238,https://old.reddit.com/r/Jokes/comments/4pqcp0/the_2016_nba_draft/,self.jokes,,[deleted],The 2016 NBA draft...,0
post,4pqcah,2qh72,jokes,false,1466818076,https://old.reddit.com/r/Jokes/comments/4pqcah/when_trump_and_boris_are_elected/,self.jokes,,"&gt;When Trump and Boris are elected...

...they'll be like toupees in a pod.",When Trump and Boris are elected...,2
post,4pqb1j,2qh72,jokes,false,1466817529,https://old.reddit.com/r/Jokes/comments/4pqb1j/why_did_princess_diana_cross_the_road/,self.jokes,,[deleted],Why did princess Diana cross the road?,0
post,4pqayu,2qh72,jokes,false,1466817488,https://old.reddit.com/r/Jokes/comments/4pqayu/how_much_space_is_left_in_the_eu/,self.jokes,,[removed],How much space is left in the EU?,2
post,4pqaol,2qh72,jokes,false,1466817374,https://old.reddit.com/r/Jokes/comments/4pqaol/the_european_union/,self.jokes,,[deleted],The European Union,1
post,4pqao3,2qh72,jokes,false,1466817368,https://old.reddit.com/r/Jokes/comments/4pqao3/did_you_hear_about_the_irish_ice_factory/,self.jokes,,They now export to Britain since the Brits thought the recipe was an EU regulation.,Did you hear about the Irish ice factory?,0
post,4pqab3,2qh72,jokes,false,1466817197,https://old.reddit.com/r/Jokes/comments/4pqab3/what_did_the_traffic_light_say_to_the_other/,self.jokes,,Don't look i'm changing,what did the traffic light say to the other traffic light?,2
post,4pqa4g,2qh72,jokes,false,1466817110,https://old.reddit.com/r/Jokes/comments/4pqa4g/what_does_britain_and_a_young_catholic_couple/,self.jokes,,[deleted],What does Britain and a young catholic couple have in common?,0
post,4pqa3r,2qh72,jokes,false,1466817102,https://old.reddit.com/r/Jokes/comments/4pqa3r/there_are_so_many_pakistanis_and_nigerians_in/,self.jokes,,The city is starting to feel a lot less Polish,There are so many Pakistanis and Nigerians in London these days,1
post,4pq9zz,2qh72,jokes,false,1466817053,https://old.reddit.com/r/Jokes/comments/4pq9zz/tifu/,self.jokes,,By posting a really stupid joke on reddit. ,TIFU....,0
post,4pq9yg,2qh72,jokes,false,1466817039,https://old.reddit.com/r/Jokes/comments/4pq9yg/i_dont_want_to_bash_jews/,self.jokes,,but come on for christ's sake.  They're bad people.,I don't want to bash jews,0
post,4pq9nr,2qh72,jokes,false,1466816903,https://old.reddit.com/r/Jokes/comments/4pq9nr/who_did_the_philosophy_major_ask_out_for_the/,self.jokes,,Nobody. He was too 'Freud. ,Who did the philosophy major ask out for the Halloween dance?,0
post,4pq9bp,2qh72,jokes,false,1466816761,https://old.reddit.com/r/Jokes/comments/4pq9bp/ive_consulted_with_my_wife/,self.jokes,,[deleted],Ive consulted with my wife..,1
post,4pq9a7,2qh72,jokes,false,1466816740,https://old.reddit.com/r/Jokes/comments/4pq9a7/a_man_comes_home_and_tells_his_wife_honey_were/,self.jokes,,"She says ""No, I hate hunting!"" 

He says ""either we're going hunting, or I'm fucking you in the ass AND you're giving me a blowjob""

The wife replies ""Alright listen, I'm not going hunting, and I'm not gonna let you fuck me in the ass, but I'll give you a blowjob"" He begrudgingly agrees. When she unzips his pants a horrible smell comes out. She takes one whiff and backs away, asking ""Honey your dick... it smells so bad, I can't go down on you... what is that?""

He angrily zips up his pants and replies ""Yeah well the dogs didn't wanna go hunting either.""
","A man comes home and tells his wife ""Honey, we're going hunting!""",16
post,4pq93n,2qh72,jokes,false,1466816651,https://old.reddit.com/r/Jokes/comments/4pq93n/with_the_way_the_value_of_the_pound_took_a/,self.jokes,,"... Instead of Brexit, they should have called it the Great Brecession.",With the way the value of the pound took a nosedive today...,2
post,4pq91b,2qh72,jokes,false,1466816623,https://old.reddit.com/r/Jokes/comments/4pq91b/i_ate_four_bowls_of_alphabet_soup/,self.jokes,,Then I had a massive vowel movement,I ate four bowls of Alphabet Soup...,110
post,4pq8z8,2qh72,jokes,false,1466816600,https://old.reddit.com/r/Jokes/comments/4pq8z8/what_kind_of_glass_do_they_put_up_in_restaurant/,self.jokes,,Hunger panes.,What kind of glass do they put up in restaurant windows to make people want to eat more?,2
post,4pq8r1,2qh72,jokes,false,1466816501,https://old.reddit.com/r/Jokes/comments/4pq8r1/what_do_you_call_a_ghost_turd/,self.jokes,,[deleted],What do you call a ghost turd?,35
post,4pq8gp,2qh72,jokes,false,1466816368,https://old.reddit.com/r/Jokes/comments/4pq8gp/now_that_brexit_is_over/,self.jokes,,"we can expect 

1. Nexit
2. Frexit 
3. Grexit 
4. Departugal 
5. Italeave
6. Czechout
7. Outstria 
8. Finish
9. Slovakout
10. Latervia
11. Byegium
12. Polend 
",Now that Brexit is over,6
post,4pq8f9,2qh72,jokes,false,1466816348,https://old.reddit.com/r/Jokes/comments/4pq8f9/what_do_you_call_someone_who_only_speaks_one/,self.jokes,,American,What do you call someone who only speaks one language?,1
post,4pq89a,2qh72,jokes,false,1466816284,https://old.reddit.com/r/Jokes/comments/4pq89a/my_girl_says_im_like_a_volcano_in_bed/,self.jokes,,Dormant,My girl says I'm like a volcano in bed...,15
post,4pq7z7,2qh72,jokes,false,1466816164,https://old.reddit.com/r/Jokes/comments/4pq7z7/why_are_pills_white/,self.jokes,,Because they work.,Why are pills white?,9
post,4pq7vw,2qh72,jokes,false,1466816118,https://old.reddit.com/r/Jokes/comments/4pq7vw/did_you_hear_how_canada_got_its_name/,self.jokes,,"The leaders couldn't decide on a name for their nation so they decided to grab a scrabble bag and choose 3 random letters.

One of the leaders sticks his hand into the bag and picks a letter out.   He then announces the letter to the leaders.

""C...ay""

Goes for the next letter and announces that.  ""N...ay"".

Finally goes for one more letter.  ""D...ay""

Edit: told it twice on accident.",Did you hear how Canada got its name?,1
post,4pq7ph,2qh72,jokes,false,1466816048,https://old.reddit.com/r/Jokes/comments/4pq7ph/did_you_know_a_cat_can_jump_higher_than_a_house/,self.jokes,,This is due to the fact that cats have very powerful hind legs and that houses can't jump.,Did you know a cat can jump higher than a house?,45
post,4pq7js,2qh72,jokes,false,1466815973,https://old.reddit.com/r/Jokes/comments/4pq7js/the_old_rooster/,self.jokes,,"An old farmer decided it was time to get a new rooster for his hens. The current rooster was still doing an okay job, but he was getting on in years and the farmer figured getting a new rooster couldn't hurt. So he buys a new cock from the local rooster emporium, and turns him loose in the barnyard. Well, the old rooster sees the young one strutting around and he's a little worried about being replaced. He walks up to the new bird.
""So you're the new stud in town? I bet you really think you're hot stuff don't you? Well I'm not ready for the chopping block yet. I'll bet I'm still the better bird. And to prove it, I challenge you to a race around that hen house over there. We'll run around it ten times and whoever finishes first gets to have all the hens for himself.""
Well, the young rooster was a proud sort, and he definitely thought he was more than a match for the old guy.
""You're on,"" he said, ""and since I'm so great, I'll even give you a head start of half a lap. I'll still win easy!""
So the two roosters go over to the henhouse to start the race with all the hens gathering to watch. The race begins and all the hens start cheering the old rooster on. After the first lap, the old rooster is still maintaining his lead.
After the second lap, the old guy's lead has slipped a little -- but he's still hanging in there. Unfortunately, the old rooster's lead continues to slip each time around, and by the fifth lap he's just barely in front of the young fella. By now the farmer has heard the commotion. He runs into the house, gets his shotgun and runs into the barnyard figuring a fox or something is after his chickens. When he gets there, he sees the two roosters running around the hen house, with the old rooster still slightly in the lead. He immediately takes his shotgun, aims, fires, and blows the young rooster away.
""Damn. That's the third gay rooster I've bought this month.""",The old rooster.,3
post,4pq7ha,2qh72,jokes,false,1466815940,https://old.reddit.com/r/Jokes/comments/4pq7ha/the_pound/,self.jokes,,[removed],The pound,1
post,4pq6p1,2qh72,jokes,false,1466815603,https://old.reddit.com/r/Jokes/comments/4pq6p1/afraid/,self.jokes,,Alone in my room and and thinking someone is also there lol.,afraid,0
post,4pq6l3,2qh72,jokes,false,1466815551,https://old.reddit.com/r/Jokes/comments/4pq6l3/a_man_who_feels_like_a_woman_consults_a_doctor/,self.jokes,,[deleted],A man who feels like a woman consults a doctor.,0
post,4pq6d9,2qh72,jokes,false,1466815460,https://old.reddit.com/r/Jokes/comments/4pq6d9/im_really_obsessed_with_harry_potter_on_a_scale/,self.jokes,,9 3/4,"I'm really obsessed with Harry Potter. On a scale of 1-10, how obsessed do you think I am?",0
post,4pq640,2qh72,jokes,false,1466815355,https://old.reddit.com/r/Jokes/comments/4pq640/whats_an_fbi_agents_favorite_feature_on_youtube/,self.jokes,,The watchlist.,What's an FBI agent's favorite feature on YouTube?,3
post,4pq62q,2qh72,jokes,false,1466815340,https://old.reddit.com/r/Jokes/comments/4pq62q/what_do_you_call_a_bear_that_is_not_jewish/,self.jokes,,Gentile Ben,What do you call a bear that is not Jewish?,3
post,4pq5tt,2qh72,jokes,false,1466815240,https://old.reddit.com/r/Jokes/comments/4pq5tt/my_friend_said_the_creator_of_spiderman_took_a/,self.jokes,,He apparently called it a Stan Lee Steamer,My friend said the creator of Spider-Man took a crap on he chest.,0
post,4pq5pl,2qh72,jokes,false,1466815188,https://old.reddit.com/r/Jokes/comments/4pq5pl/can_someone_explain_that_brexit_joke/,self.jokes,,[deleted],Can someone explain that brexit joke,0
post,4pq5no,2qh72,jokes,false,1466815170,https://old.reddit.com/r/Jokes/comments/4pq5no/i_used_to_be_fat/,self.jokes,,[deleted],I used to be fat,0
post,4pq5bn,2qh72,jokes,false,1466815041,https://old.reddit.com/r/Jokes/comments/4pq5bn/just_went_to_my_local_asda_tonight/,self.jokes,,"Just been to my local Asda and there was a Polish couple in front of me, the cashier asked do you want help packing your bags? 

I thought bloody hell this is happening faster than I thought!",Just went to my local asda tonight...,1
post,4pq4cr,2qh72,jokes,false,1466814670,https://old.reddit.com/r/Jokes/comments/4pq4cr/how_can_you_spot_a_blind_guy_at_a_nudist_colony/,self.jokes,,It's not hard.,How can you spot a blind guy at a nudist colony?,2
post,4pq4bv,2qh72,jokes,false,1466814659,https://old.reddit.com/r/Jokes/comments/4pq4bv/brexit/,self.jokes,,EU now has 1 GB of free space!!,Brexit,0
post,4pq417,2qh72,jokes,false,1466814539,https://old.reddit.com/r/Jokes/comments/4pq417/jk_rowling_hid_some_text_on_the_title_of_harry/,self.jokes,,[deleted],J.K. Rowling hid some text on the title of Harry Potter,0
post,4pq2nb,2qh72,jokes,false,1466813956,https://old.reddit.com/r/Jokes/comments/4pq2nb/two_jewish_guys_walking_down_the_street_see_a/,self.jokes,,[deleted],"Two Jewish guys walking down the street see a sign that says ""Christian conversions: $20.""",0
post,4pq2aw,2qh72,jokes,false,1466813825,https://old.reddit.com/r/Jokes/comments/4pq2aw/the_british_pound_has_been_given_a_new_name_to/,self.jokes,,It's called Britcoin.,The British pound has been given a new name to better represent its future stability.,1
post,4pq0qx,2qh72,jokes,false,1466813214,https://old.reddit.com/r/Jokes/comments/4pq0qx/im_not_really_that_surprised_that_there_was_a/,self.jokes,,"After all, she *is* an offensive hero.",I'm not really that surprised that there was a controversy over that Tracer pose in Overwatch.,2
post,4pq0jf,2qh72,jokes,false,1466813128,https://old.reddit.com/r/Jokes/comments/4pq0jf/whats_the_difference_between_a_feminist_and_a/,self.jokes,,A spear has a point,What's the difference between a feminist and a spear...,8
post,4pq0e9,2qh72,jokes,false,1466813075,https://old.reddit.com/r/Jokes/comments/4pq0e9/two_of_my_favourite_moments_in_my_life_were_when/,self.jokes,,I hit him so hard he slept through the whole thing,Two of my favourite moments in my life were when I won my first fight and lost my virginity,11
post,4pq078,2qh72,jokes,false,1466813000,https://old.reddit.com/r/Jokes/comments/4pq078/there_was_a_girl_who_went_to_a_park/,self.jokes,,[deleted],There was a girl who went to a park,0
post,4pq03u,2qh72,jokes,false,1466812964,https://old.reddit.com/r/Jokes/comments/4pq03u/i_guess_the_eu/,self.jokes,,[deleted],I guess the EU ...,0
post,4pq029,2qh72,jokes,false,1466812945,https://old.reddit.com/r/Jokes/comments/4pq029/what_does_the_doctor_say_after_colonoscopy/,self.jokes,,"See ewwww later!
",What does the doctor say after colonoscopy?,0
post,4ppzq5,2qh72,jokes,false,1466812804,https://old.reddit.com/r/Jokes/comments/4ppzq5/france_to_britain_after_the_brexit_vote_leave/,self.jokes,,[removed],"France to Britain after the Brexit vote: ""Leave right away, and good riddance, we've never needed you for anything ever anyhow""",1
post,4ppzpo,2qh72,jokes,false,1466812800,https://old.reddit.com/r/Jokes/comments/4ppzpo/whats_the_difference_between_a_chickpea_and_a/,self.jokes,,...I've never had a garbanzo bean on my face,What's the difference between a chickpea and a garbanzo bean?,1
post,4ppzfl,2qh72,jokes,false,1466812693,https://old.reddit.com/r/Jokes/comments/4ppzfl/i_wonder_what_the_first_holocaust_joke_ever_made/,self.jokes,,[deleted],I wonder what the first Holocaust joke ever made was...,0
post,4ppzey,2qh72,jokes,false,1466812688,https://old.reddit.com/r/Jokes/comments/4ppzey/never_knew_that_irish_people_are_so_racist/,self.jokes,,Needless to say I was shocked when my Irish mate started telling me about how much he hates the black and tans.,Never knew that Irish people are so racist...,1
post,4ppzdj,2qh72,jokes,false,1466812670,https://old.reddit.com/r/Jokes/comments/4ppzdj/i_heard_somewhere_that/,self.jokes,,"You only remember things that you read, is that true?",I heard somewhere that...,0
post,4ppz3k,2qh72,jokes,false,1466812555,https://old.reddit.com/r/Jokes/comments/4ppz3k/you_gotta_hand_it_to_leave_brits/,self.jokes,,They were so concerned about immigrants ruining their economy that they preempted it and ruined their economy themselves.,You Gotta Hand It To Leave Brits,0
post,4ppz1t,2qh72,jokes,false,1466812532,https://old.reddit.com/r/Jokes/comments/4ppz1t/a_muslim_walks_into_a_bar_and_says/,self.jokes,,[removed],a muslim walks into a bar and says,1
post,4ppyvf,2qh72,jokes,false,1466812457,https://old.reddit.com/r/Jokes/comments/4ppyvf/an_atheist_a_vegan_and_a_crossfitter_walk_into_a/,self.jokes,,[deleted],"An atheist, a vegan, and a crossfitter walk into a bar...",0
post,4ppyjk,2qh72,jokes,false,1466812315,https://old.reddit.com/r/Jokes/comments/4ppyjk/what_does_the_doctor_say_after_colonoscopy/,self.jokes,,[deleted],What does the doctor say after colonoscopy?,0
post,4ppydp,2qh72,jokes,false,1466812241,https://old.reddit.com/r/Jokes/comments/4ppydp/i_guess_the_eu/,self.jokes,,[deleted],I guess the EU ...,1
post,4ppy6t,2qh72,jokes,false,1466812172,https://old.reddit.com/r/Jokes/comments/4ppy6t/in_tesco_earlier/,self.jokes,,"the cashier asked the Foreign couple in front of me if they wanted help packing their bags. Fuck me, we only voted out yesterday, give them a chance!!!",In Tesco earlier,2
post,4ppxuz,2qh72,jokes,false,1466812032,https://old.reddit.com/r/Jokes/comments/4ppxuz/i_stopped_feeling_empty_inside_today_after_a_long/,self.jokes,,But then I pooped,I stopped feeling empty inside today after a long fight with anxiety/depression.,0
post,4ppxda,2qh72,jokes,false,1466811827,https://old.reddit.com/r/Jokes/comments/4ppxda/the_five_senses_are_touch_smell_sight_hearing_and/,self.jokes,,It's on the tip of my tongue...,"The five senses are touch, smell, sight, hearing, and.....",6
post,4ppwts,2qh72,jokes,false,1466811630,https://old.reddit.com/r/Jokes/comments/4ppwts/two_men_from_texas_were_sitting_at_a_bar/,self.jokes,,"Two men from Texas were sitting at a bar, when a young lady nearby began to choke on a hamburger. She gasped and gagged, and one Texan turned to the other and said, ""That little gal is havin' a bad time. I'm a gonna go over there and help."" He ran over to the young lady, held both sides of her head in his big, Texan hands, and asked, ""Kin ya swaller?"" Gasping, she shook her head no. He asked, ""Kin ya breathe?"" Still gasping, she again shook her head no. With that, he yanked up her skirt, pulled down her panties and licked her on the butt. The young woman was so shocked that she coughed up the piece of hamburger and began to breathe on her own. The Texan sat back down with his friend and said, ""Ya know, it's sure amazin' how that hind-lick manoeuvre always works.""",Two men from Texas were sitting at a bar,23
post,4ppwq6,2qh72,jokes,false,1466811590,https://old.reddit.com/r/Jokes/comments/4ppwq6/a_joke_for_dumb_people/,self.jokes,,"okay dont kill me just yet lol okay 
okay a Jewish mom goes soccer league in Ireland and she says ""excuse me sir do you know where i can get a soccer player from?"" then the irish man says ""no ma'am you dont buy them you watch them play fut ball"" and the jewish mom says ""well my irene i need to kidnap one then and make them my husband"" then an soccer player comes up to her and gives her a beer and makes her play soccer. an hour later she got on the soccer team and every time she would play she would always drink the blood of germans",a joke for dumb people,0
post,4ppw2w,2qh72,jokes,false,1466811337,https://old.reddit.com/r/Jokes/comments/4ppw2w/great_britain_is_leaving_the_eu/,self.jokes,,"Markets are panicked.  Countries are worried.  N. Ireland and Scotland may leave, leaving Great Britain as just Britain.

What would they call the new land of N. Ireland and Scotland?  Great Scott!",Great Britain is leaving the EU,0
post,4ppvve,2qh72,jokes,false,1466811247,https://old.reddit.com/r/Jokes/comments/4ppvve/i_have_a_pill_that_helps_you_lose_pounds_fast/,self.jokes,,its called the brexit pill,I have a pill that helps you lose pounds fast,0
post,4ppvov,2qh72,jokes,false,1466811174,https://old.reddit.com/r/Jokes/comments/4ppvov/did_you_know_that_all_milk_has_to_be_sterilized/,self.jokes,,Prepasteurous!,Did you know that all milk has to be sterilized before use?,6
post,4ppvoq,2qh72,jokes,false,1466811172,https://old.reddit.com/r/Jokes/comments/4ppvoq/i_guess_the_eu_has_1_gb_of_free_space_now/,self.jokes,,[removed],I guess the EU has 1 GB of free space now...,1
post,4ppv7p,2qh72,jokes,false,1466810978,https://old.reddit.com/r/Jokes/comments/4ppv7p/a_group_of_jews_went_to_auschwitz_for_vacation/,self.jokes,,"They gave it one star.
",A Group of Jews went to Auschwitz for Vacation,0
post,4ppumy,2qh72,jokes,false,1466810749,https://old.reddit.com/r/Jokes/comments/4ppumy/where_do_most_pirates_come_from/,self.jokes,,Arrrrgentina,Where do most pirates come from?,0
post,4ppumi,2qh72,jokes,false,1466810745,https://old.reddit.com/r/Jokes/comments/4ppumi/you_know_you_might_be_a_prison_officer_when/,self.jokes,,"1. You have the bladder capacity of five people.
2. You have ever restrained someone and it was not a sexual experience.
3. You believe at least 50% of people are a waste of skin.
4. Your idea of a good time is a cell entry at shift change.
5. You do a strip search on anyone who seems remotely friendly towards you.
6. Discussing dismemberment over a gourmet meal seems perfectly normal.
7. You find humour in other people's stupidity.
8. You believe in aerial spraying of Prozac.
9. Your idea of comforting an prisoner is placing him in full bed restraints.
10. You believe that ""shallow gene pool"" is sufficient grounds for a misconduct report.
11. You believe the government should require extensive testing and permits prior to reproduction.
12. You believe that unspeakable evils will befall you if anyone says ""Boy, it sure is quiet around here.""
13. Your diet consists of food that has gone through more processing than a computer can track.
14. You believe chocolate is a food group.
15. You have contemplated holding a seminar titled ""SUICIDE - Getting It Right The First Time.""
16. You believe that ""Too stupid to live"" is a valid verdict.
17. You have to put the phone down before you begin laughing uncontrollably.
18. You think caffeine should be available in IV form.
19. Your favourite hallucinogen is exhaustion.
20. When you mention ""vegetables,"" you are not referring to the food group.
21. It occurs to you one night that you really have entered, ""The Twilight Zone.""
22. You find out a lot about paranoia just by following prisoners around.
23. You're escorting a smurf to clinical and find yourself carrying on an intelligent conversation with him.
24. You believe it's not a good riot unless it involves overtime.
25. You are the only person introduced by profession at a social gathering.
26. You walk into places and people think it highly comical to seize a co-worker and shout, ""They've come to get you Frank!""
27. People shout, ""I didn't do it!"" when you walk into the room in uniform and they think they are being hysterically funny and original.
28. You believe in involuntary sterilization.
29. You had to work 18 years to earn what the rookies are starting at now.
30. When you mention ""Bugs"", you are not referring to insects.
",You know you might be a Prison Officer when:,0
post,4ppu4x,2qh72,jokes,false,1466810557,https://old.reddit.com/r/Jokes/comments/4ppu4x/i_guess_eu_has_1_gb_of_free_space_now/,self.jokes,,[removed],I guess EU has 1 GB of free space now...,1
post,4pptvj,2qh72,jokes,false,1466810458,https://old.reddit.com/r/Jokes/comments/4pptvj/a_political_joke_for_americans/,self.jokes,,I'm voting for hillary,A political joke for Americans,0
post,4pptql,2qh72,jokes,false,1466810397,https://old.reddit.com/r/Jokes/comments/4pptql/what_is_the_easiest_way_to_know_if_a_rabbit_is/,self.jokes,,His carrot smells like shit,What is the easiest way to know if a rabbit is homosexual?,6
post,4ppsvs,2qh72,jokes,false,1466810048,https://old.reddit.com/r/Jokes/comments/4ppsvs/whats_the_difference_between_a_sociopath_and_a/,self.jokes,,You can't ride your bike on a sociopath,What's the difference between a sociopath and a psychopath?,4
post,4ppsg6,2qh72,jokes,false,1466809868,https://old.reddit.com/r/Jokes/comments/4ppsg6/what_did_gb_say_to_eu/,self.jokes,,"Peace out, EUROn EUROwn!",What did GB say to EU?,7
post,4ppsez,2qh72,jokes,false,1466809854,https://old.reddit.com/r/Jokes/comments/4ppsez/one_night_as_a_couple_lay_down_to_bed/,self.jokes,,"the husband gently starts rubbing his wife on the arm. The wife turned over and said ""Sorry honey, I have an OBGYN appointment tomorrow and I want to stay fresh.""

Dejected and rejected, the hubby tries to sleep. After a while he turns over to his wife and says ""Do you have a dentist's appointment too?""
","One Night, as a couple lay down to bed,",14
post,4pps4a,2qh72,jokes,false,1466809739,https://old.reddit.com/r/Jokes/comments/4pps4a/tifu_by_eating_my_coworkers_sandwich/,self.jokes,,"Oops, wrong sub",TIFU by eating my coworkers sandwich,18
post,4pps32,2qh72,jokes,false,1466809731,https://old.reddit.com/r/Jokes/comments/4pps32/whats_2_blink_182/,self.jokes,,46,What's 2 + Blink 182,2
post,4pprw6,2qh72,jokes,false,1466809659,https://old.reddit.com/r/Jokes/comments/4pprw6/what_happens_when_david_cameron_gets_a_gift/,self.jokes,,[deleted],What happens when David Cameron gets a gift basket he isn't pleased with?,1
post,4ppr8n,2qh72,jokes,false,1466809418,https://old.reddit.com/r/Jokes/comments/4ppr8n/insomnia_is_very_common/,self.jokes,,Try not to lose any sleep over it.,Insomnia is very common.,24
post,4ppr7v,2qh72,jokes,false,1466809412,https://old.reddit.com/r/Jokes/comments/4ppr7v/son_in_college_sends_his_dad_a_text/,self.jokes,,[removed],Son in college sends his dad a text...,1
post,4ppqmz,2qh72,jokes,false,1466809208,https://old.reddit.com/r/Jokes/comments/4ppqmz/whats_the_great_way_to_lose_some_pounds/,self.jokes,,Leave the EU.,Whats the great way to lose some pounds?,0
post,4ppqia,2qh72,jokes,false,1466809151,https://old.reddit.com/r/Jokes/comments/4ppqia/whats_the_difference_between_a_pound_and_a_dollar/,self.jokes,,A dollar,What's the difference between a Pound and a Dollar?,345
post,4pppo4,2qh72,jokes,false,1466808819,https://old.reddit.com/r/Jokes/comments/4pppo4/a_farmer_is_oppressing_his_chickens/,self.jokes,,[removed],A Farmer is Oppressing his chickens...,1
post,4pppln,2qh72,jokes,false,1466808796,https://old.reddit.com/r/Jokes/comments/4pppln/had_to_get_a_colonoscopy_today/,self.jokes,,It was a real pain the ass. ,Had to get a colonoscopy today,3
post,4pppjw,2qh72,jokes,false,1466808775,https://old.reddit.com/r/Jokes/comments/4pppjw/before_it_starts/,self.jokes,,"A man came home from work, sat down in his favourite chair, turned on the TV, and said to his wife, ""Quick, bring me a beer before it starts""

She looked a little puzzled, but brought him a beer. When he finished it, he said, ""Quick, bring me another beer. It's gonna start.""

This time she looked a little angry, but brought him a beer.

When it was gone, he said, ""Quick, another beer before it starts.""

""That's it!"" She blows her top, ""You bastard! You waltz in here, flop your fat ass down, don't even say hello to me and then expect me to run around like your slave. Don't you realize that I cook and clean and wash and iron all day long?""

The husband sighed. ""Oh shit, it started!”
",Before it starts...,115
post,4pppei,2qh72,jokes,false,1466808720,https://old.reddit.com/r/Jokes/comments/4pppei/if_france_leaves_the_eu/,self.jokes,,They would be disenfrance-ised.,If France leaves the EU....,1
post,4ppp8l,2qh72,jokes,false,1466808659,https://old.reddit.com/r/Jokes/comments/4ppp8l/a_man_is_walking_down_the_beach/,self.jokes,,"He see's a sign that says, ""$50 blow job, while singing"". 

He scratches his head and decides, what the heck. So he goes in, there is this pretty attractive woman, so he puts down his $50. She starts giving him an amazing blow job and right in the middle, she pipes up with this incredible singing voice. 

The man leaves and goes home. Later that night, he just can't figure out what's happening. So he goes back the next day and puts his $50 down. She turns off the lights, another amazing blow job and half way thru, the singing begins. It's definitely not a recording. It's her voice for sure

He leaves but can't shake the confusion. So he deduces a plan. The next day he returns and puts down his $50. She turns off the lights, once again, gives an amazing blow job and in the middle, she starts singing.

Then he reaches over, turns on the lights and there is a glass eye ball on the table. ",A man is walking down the beach,8
post,4ppoug,2qh72,jokes,false,1466808508,https://old.reddit.com/r/Jokes/comments/4ppoug/brexit_to_be_followed_by_grexit_departugal/,self.jokes,,[removed],'Brexit' to be followed by Grexit. Departugal. Italeave. Fruckoff. Czechout. Oustria. Finish. Slovakout. Latervia. Byegium.,1
post,4ppnyh,2qh72,jokes,false,1466808168,https://old.reddit.com/r/Jokes/comments/4ppnyh/what_do_you_purchase_paintings_with/,self.jokes,,[removed],What do you purchase paintings with?,1
post,4ppnwf,2qh72,jokes,false,1466808151,https://old.reddit.com/r/Jokes/comments/4ppnwf/what_have_disney_and_the_uk_got_in_common/,self.jokes,,Both dropped the EU And screwed over a lot of people,What have Disney and the U.K. got in common?,4
post,4ppnps,2qh72,jokes,false,1466808081,https://old.reddit.com/r/Jokes/comments/4ppnps/hope_you_enjoy_it/,self.jokes,,Why do women live on average two years longer? Because the time they spend parking doesn’t count.,Hope you enjoy it,5
post,4ppnis,2qh72,jokes,false,1466808000,https://old.reddit.com/r/Jokes/comments/4ppnis/what_did_paul_revere_say_last_night/,self.jokes,,"The British are coming, the British are coming!",What did Paul Revere say last night?,0
post,4ppmv4,2qh72,jokes,false,1466807749,https://old.reddit.com/r/Jokes/comments/4ppmv4/whats_the_difference_between_bill_clinton_and/,self.jokes,,Hillary won't suck Bill's dick.,What's the difference between Bill Clinton and Israel?,5
post,4ppmm0,2qh72,jokes,false,1466807656,https://old.reddit.com/r/Jokes/comments/4ppmm0/hello_how_many_british_persons_does_it_take_to/,self.jokes,,I'll tell you. One to screw in the lightbulb and sixty-four million to vote on a referendum about whether or not to stay in the dark. ,Hello. How many British persons does it take to change a lightbulb?,0
post,4ppm91,2qh72,jokes,false,1466807521,https://old.reddit.com/r/Jokes/comments/4ppm91/to_all_those_people_that_have_ever_talked_about/,self.jokes,,You discussed me.,To all those people that have ever talked about me behind my back...,7
post,4ppm34,2qh72,jokes,false,1466807452,https://old.reddit.com/r/Jokes/comments/4ppm34/snoop_and_dre_might_be_getting_old_but_at_least/,self.jokes,,"Their new album is called ""Pissin' Aint Easy, But Its Necessary"".   ","Snoop and Dre might be getting old, but at least they still keeping it real..",0
post,4pplwz,2qh72,jokes,false,1466807396,https://old.reddit.com/r/Jokes/comments/4pplwz/why_do_all_women_like_jesus/,self.jokes,,[deleted],Why do all women like Jesus?,1
post,4ppluo,2qh72,jokes,false,1466807377,https://old.reddit.com/r/Jokes/comments/4ppluo/theres_now_more_free_space_in_the_european_union/,self.jokes,,[deleted],There's now more free space in the European Union,1
post,4pplsn,2qh72,jokes,false,1466807359,https://old.reddit.com/r/Jokes/comments/4pplsn/george_went_on_a_vacation_to_the_middle_east/,self.jokes,,"George went on a vacation to the Middle East with most of his family, including his mother-in-law.  During their vacation, and while they were visiting Jerusalem, George's mother-in-law died.  With the death certificate in hand, George went to the American Consulate Office to make arrangements to send the body back to the States for proper burial.  The Consul, after hearing of the death of the mother-in-law, told George, 

""My friend, the sending of a body back to the States for burial is very, very expensive.  It could cost as much as $5,000 dollars.""  The Consul continued, ""In most of these cases, the person responsible for the remains normally decides to bury the body here.  This would only cost $150 dollars"".  

George thinks for some time, and answers the Consul, 

""I don't care how much it will cost to send the body back.  That's what I want to do.""  

The Consul, after hearing this says, ""You must have loved your mother-in-law very much, considering the difference in price between $5,000 and $150 dollars.""  

""No, it's not that,"" says George.  ""You see, I know of a case many, many years ago of a person that was buried here in Jerusalem, and on the third day he was resurrected.  Consequently, I do not want to take that chance!""
",George went on a vacation to the Middle East...,21
post,4ppleb,2qh72,jokes,false,1466807216,https://old.reddit.com/r/Jokes/comments/4ppleb/an_old_woman_and_her_poolboy/,self.jokes,,"An old woman catches her long time poolboy rummaging through her drawers one day.
""Pervert!"" She screams. ""You will be punished for this!""
""Now, take off my shoes""
And the poolboy takes off her shoes.
""Now my stockings.""
He takes off her stockings.
""Now unbutton my blouse!"" 
He does, reluctantly.
""And lastly, my bra.""
The poolboy weeps as he does what he's told.
The old woman looks at him sternly and says....

""If I EVER catch you wearing my clothes again, you're fired!""",An old woman and her poolboy...,0
post,4ppl9c,2qh72,jokes,false,1466807177,https://old.reddit.com/r/Jokes/comments/4ppl9c/do_you_know_what_would_a_genetic_crossover/,self.jokes,,[deleted],Do you know what would a genetic crossover between a black man and an octopus look like?,0
post,4ppkaq,2qh72,jokes,false,1466806821,https://old.reddit.com/r/Jokes/comments/4ppkaq/im_a_little_late_with_the_uk_leaving_the_eu_news/,self.jokes,,[deleted],Im a little late with the UK leaving the EU news,0
post,4ppk0a,2qh72,jokes,false,1466806714,https://old.reddit.com/r/Jokes/comments/4ppk0a/so_how_we_call_uk_after_brexit/,self.jokes,,[deleted],So how we call UK after Brexit?,0
post,4ppjyv,2qh72,jokes,false,1466806697,https://old.reddit.com/r/Jokes/comments/4ppjyv/why_was_it_hard_to_talk_to_polish_people_in_1938/,self.jokes,,[deleted],Why was it hard to talk to Polish people in 1938?,1
post,4ppjrv,2qh72,jokes,false,1466806627,https://old.reddit.com/r/Jokes/comments/4ppjrv/a_muslim_who_isnt_a_terrorist/,self.jokes,,[removed],A Muslim who isn't a terrorist...,1
post,4ppjph,2qh72,jokes,false,1466806602,https://old.reddit.com/r/Jokes/comments/4ppjph/when_donald_trump_wins_the_election_the_top/,self.jokes,,[removed],"When Donald Trump wins the election, the top Google search result for voters in the U.S. will be ""How to commit 'sudoku'""",1
post,4ppjnc,2qh72,jokes,false,1466806581,https://old.reddit.com/r/Jokes/comments/4ppjnc/scotland_highly_likely_to_have_another/,self.jokes,,[deleted],Scotland highly likely to have another independence referendum,3
post,4ppjj9,2qh72,jokes,false,1466806542,https://old.reddit.com/r/Jokes/comments/4ppjj9/whats_another_name_for_a_teepee/,self.jokes,,Injinuity,What's another name for a teepee?,0
post,4ppitq,2qh72,jokes,false,1466806273,https://old.reddit.com/r/Jokes/comments/4ppitq/what_do_you_call_batman_when_he_skips_church/,self.jokes,,[deleted],What do you call Batman when he skips church?,0
post,4ppi1t,2qh72,jokes,false,1466805994,https://old.reddit.com/r/Jokes/comments/4ppi1t/if_i_had_100_pounds/,self.jokes,,[deleted],If i had 100 pounds...,0
post,4pphp2,2qh72,jokes,false,1466805869,https://old.reddit.com/r/Jokes/comments/4pphp2/a_muslim_man_sends_his_son_to_mecca/,self.jokes,,[deleted],A Muslim man sends his son to Mecca ...,0
post,4ppgc1,2qh72,jokes,false,1466805356,https://old.reddit.com/r/Jokes/comments/4ppgc1/joke/,self.jokes,,"Police officer: ""Can you identify yourself, sir?""
 
Driver pulls out his mirror and says: ""Yes, it's me.""",Joke,15
post,4ppfv8,2qh72,jokes,false,1466805183,https://old.reddit.com/r/Jokes/comments/4ppfv8/trump_to_britain/,self.jokes,,[deleted],Trump to Britain......,2
post,4ppfsg,2qh72,jokes,false,1466805157,https://old.reddit.com/r/Jokes/comments/4ppfsg/want_to_lose_some_weight_well_head_over_to_great/,self.jokes,,"Want to lose some weight? Too tired always running on the treadmill? Well we've got the solution for you. Head on over to Great Britain, you'll drop some quick pounds.",Want to lose some weight? Well head over to Great Britain.,0
post,4ppfp7,2qh72,jokes,false,1466805123,https://old.reddit.com/r/Jokes/comments/4ppfp7/what_does_david_cameron_and_a_one_night_stand/,self.jokes,,[deleted],What does David Cameron and a one night stand have in common?,3
post,4ppfdn,2qh72,jokes,false,1466805013,https://old.reddit.com/r/Jokes/comments/4ppfdn/i_just_asked_my_dad_what_his_favourite_part_about/,self.jokes,,"He responded with June, July, and August",I just asked my dad what his favourite part about being a teacher is...,9
post,4ppetd,2qh72,jokes,false,1466804814,https://old.reddit.com/r/Jokes/comments/4ppetd/what_does_a_mexican_duck_say/,self.jokes,,Guac guac,What does a Mexican duck say?,11
post,4ppdy1,2qh72,jokes,false,1466804495,https://old.reddit.com/r/Jokes/comments/4ppdy1/since_the_pound_has_lost_so_much_value/,self.jokes,,...maybe it should be renamed to the Ounce,Since the Pound has lost so much value...,0
post,4ppdvm,2qh72,jokes,false,1466804470,https://old.reddit.com/r/Jokes/comments/4ppdvm/redditors_of_mississippi_tell_me_how_do_you_feel/,self.jokes,,"Oh wait, you can't read.",Redditors of Mississippi. Tell me how do you feel abou-,0
post,4ppdli,2qh72,jokes,false,1466804370,https://old.reddit.com/r/Jokes/comments/4ppdli/why_does_it_cost_a_wizard_so_much_money_to_spy_on/,self.jokes,,"Well because it's ex-pensieve, of course!",Why does it cost a Wizard so much money to spy on the thoughts of his or her past girlfriend/boyfriend?,0
post,4ppcmr,2qh72,jokes,false,1466804022,https://old.reddit.com/r/Jokes/comments/4ppcmr/so_my_wife_came_up_to_me_and_said_take_off_my/,self.jokes,,"So I took off her shirt. Then she said, ""Take off my skirt."" I took off her skirt. ""Take off my shoes."" I took off her shoes. ""Now my hose, bra, and panties."" I took them off. Then she looked at me and said, ""I don't want to catch you wearing my things ever again.""","So my wife came up to me and said, ""Take off my shirt.""",0
post,4ppccv,2qh72,jokes,false,1466803926,https://old.reddit.com/r/Jokes/comments/4ppccv/whats_that_diving_is_it_a_bird_is_it_a_plane/,self.jokes,,No it's the British Pound...,"What's that diving? Is it a bird, Is it a plane...",7
post,4ppca4,2qh72,jokes,false,1466803902,https://old.reddit.com/r/Jokes/comments/4ppca4/i_have_this_great_highlighterits_called_oily_skin/,self.jokes,,i have this great highlighter its called oily skin,i have this great highlighter..its called oily skin,0
post,4ppc8p,2qh72,jokes,false,1466803888,https://old.reddit.com/r/Jokes/comments/4ppc8p/since_the_pund_has_lost_so_much_value/,self.jokes,,[deleted],Since the pund has lost so much value...,1
post,4ppc5l,2qh72,jokes,false,1466803865,https://old.reddit.com/r/Jokes/comments/4ppc5l/what_kind_of_concert_only_costs_45_cents/,self.jokes,,A British one.,What kind of concert only costs 45 cents?,0
post,4ppc1d,2qh72,jokes,false,1466803828,https://old.reddit.com/r/Jokes/comments/4ppc1d/meet_my_good_friend_50_cent_or_as_hes_known/,self.jokes,,"10,000 Pounds","Meet my good friend 50 Cent, or as he's known across the pond...",4
post,4ppbt2,2qh72,jokes,false,1466803749,https://old.reddit.com/r/Jokes/comments/4ppbt2/pork_skins_are_called_chicharones_in_spanish/,self.jokes,,I guess in China they're called chihuahuarones,Pork skins are called chicharones in Spanish...,0
post,4ppbqi,2qh72,jokes,false,1466803723,https://old.reddit.com/r/Jokes/comments/4ppbqi/australia_is_planning_to_leave_the_au/,self.jokes,,Stralia ,Australia is planning to leave the AU,0
post,4ppavd,2qh72,jokes,false,1466803403,https://old.reddit.com/r/Jokes/comments/4ppavd/did_you_hear_about_the_hooker_that_doesnt_charge/,self.jokes,,[deleted],Did you hear about the hooker that doesn't charge?,6
post,4ppasj,2qh72,jokes,false,1466803379,https://old.reddit.com/r/Jokes/comments/4ppasj/my_wife_woke_me_up_all_excited_this_morning/,self.jokes,,She said honey look at all the pounds I've lost.  I told her that she was looking at our retirement account not her fitbit.  ,My wife woke me up all excited this morning...,44
post,4ppa97,2qh72,jokes,false,1466803183,https://old.reddit.com/r/Jokes/comments/4ppa97/i_was_surprised_when_a_coworker_was_talking_about/,self.jokes,,[removed],I was surprised when a coworker was talking about the Baader-Meinhof Phenomenon. I just read about it this morning!,1
post,4ppa2f,2qh72,jokes,false,1466803119,https://old.reddit.com/r/Jokes/comments/4ppa2f/how_does_a_muslim_close_a_door/,self.jokes,,[deleted],How does a Muslim close a door?,2
post,4pp9wx,2qh72,jokes,false,1466803066,https://old.reddit.com/r/Jokes/comments/4pp9wx/try_the_brand_new_brexit_diet/,self.jokes,,[deleted],"Try the brand new ""Brexit"" diet!",0
post,4pp9u0,2qh72,jokes,false,1466803036,https://old.reddit.com/r/Jokes/comments/4pp9u0/i_regret_joining_the_gym_recently/,self.jokes,,"
Leaving the EU would've been a more effective way to lose pounds.",I regret joining the gym recently.,3
post,4pp9tx,2qh72,jokes,false,1466803034,https://old.reddit.com/r/Jokes/comments/4pp9tx/id_tell_a_corny_joke/,self.jokes,,but I'd get an earful.,I'd tell a corny joke,0
post,4pp9l5,2qh72,jokes,false,1466802943,https://old.reddit.com/r/Jokes/comments/4pp9l5/im_writing_a_fantasy_novel_like_the_works_of_jrr/,self.jokes,,[deleted],I'm writing a fantasy novel like the works of J.R.R. Tolkien.,0
post,4pp99n,2qh72,jokes,false,1466802816,https://old.reddit.com/r/Jokes/comments/4pp99n/whats_the_diving_is_it_a_bird_is_it_a_plane/,self.jokes,,[deleted],"What's the diving? Is it a bird, is it a plane...",1
post,4pp8gb,2qh72,jokes,false,1466802541,https://old.reddit.com/r/Jokes/comments/4pp8gb/two_boys_were_arguing_when_the_teacher_entered/,self.jokes,,[removed],Two boys were arguing when the teacher entered the room.,1
post,4pp89e,2qh72,jokes,false,1466802484,https://old.reddit.com/r/Jokes/comments/4pp89e/what_my_boss_just_said_today/,self.jokes,,[deleted],What my boss just said today...,1
post,4pp6y1,2qh72,jokes,false,1466802042,https://old.reddit.com/r/Jokes/comments/4pp6y1/what_do_you_call_a_black_friend/,self.jokes,,[removed],What do you call a black friend?,1
post,4pp6qb,2qh72,jokes,false,1466801965,https://old.reddit.com/r/Jokes/comments/4pp6qb/a_cop_stopped_a_man_smoking_cannabis_while_driving/,self.jokes,,"The officer asked ""how high are you?"" 
The man replied ""no officer, its hi how are you""",A cop stopped a man smoking cannabis while driving,7
post,4pp6m9,2qh72,jokes,false,1466801922,https://old.reddit.com/r/Jokes/comments/4pp6m9/i_hope_you_enjoy_this_joke/,self.jokes,,As much as my old school teacher enjoyed giving sweets to children.,I hope you enjoy this joke...,0
post,4pp6fp,2qh72,jokes,false,1466801856,https://old.reddit.com/r/Jokes/comments/4pp6fp/i_woke_up_early_today_455_am/,self.jokes,,[deleted],I woke up early today (4:55 AM),2
post,4pp5yn,2qh72,jokes,false,1466801681,https://old.reddit.com/r/Jokes/comments/4pp5yn/i_know_a_guy_who_used_to_have_leukaemia/,self.jokes,,He's Luekae to be alive.,I know a guy who used to have Leukaemia,6
post,4pp5s8,2qh72,jokes,false,1466801611,https://old.reddit.com/r/Jokes/comments/4pp5s8/the_creator_of_winrar_was_arrested_and_put_on/,self.jokes,,"The trial was supposed to last 40 days, but it keeps on going",The creator of WinRAR was arrested and put on trial,900
post,4pp5l4,2qh72,jokes,false,1466801538,https://old.reddit.com/r/Jokes/comments/4pp5l4/the_perfect_son/,self.jokes,,"The Perfect Son
A: I have the perfect son. 
B: Does he smoke? 
A: No, he doesn't. 
B: Does he drink whiskey? 
A: No, he doesn't. 
B: Does he ever come home late? 
A: No, he doesn't. 
B: I guess you really do have the perfect son. How old is he? 
A: He will be six months old next Wednesday.",The Perfect Son,0
post,4pp4tg,2qh72,jokes,false,1466801283,https://old.reddit.com/r/Jokes/comments/4pp4tg/two_jews_are_walking_down_the_street/,self.jokes,,"Moishe and Ibraham are walking down the street and they come across a church sign that says, ""Convert to Christianity! Receive $1000!"". Ibraham turns to Moishe a says, ""Well, I might as well go see what this is all about.""  
Moishe sits down on a bench and waits. He's waiting for 5 minutes, 10 minutes, an hour goes by then Ibraham finally comes out.  
Moishe says, ""So... how'd it go?""  
Ibraham replies, ""I've accepted Jesus Christ as my Lord and Savior. I believe that he died on the cross for our sins, on the third day he rose from the dead and he is now seated at the right hand of the Father.""  
Moisha says, ""What about the $1000?""  
Ibraham says, ""What is with you people and money?""  ",Two Jews are walking down the street...,222
post,4pp4k9,2qh72,jokes,false,1466801196,https://old.reddit.com/r/Jokes/comments/4pp4k9/i_woke_up_early_today/,self.jokes,,[removed],I woke up early today,1
post,4pp488,2qh72,jokes,false,1466801078,https://old.reddit.com/r/Jokes/comments/4pp488/what_do_you_call_a_kitty_thrown_out_of_a_window/,self.jokes,,[deleted],What do you call a kitty thrown out of a window?,0
post,4pp41i,2qh72,jokes,false,1466801014,https://old.reddit.com/r/Jokes/comments/4pp41i/uk_will_be_alright/,self.jokes,,[deleted],UK will be alright...,0
post,4pp3sk,2qh72,jokes,false,1466800922,https://old.reddit.com/r/Jokes/comments/4pp3sk/david_camerons_legacy/,self.jokes,,"David Cameron will go down in history as the man who fucked up his campaign, fucked up his job, and fucked up a dead pig.",David Cameron's legacy,0
post,4pp3no,2qh72,jokes,false,1466800881,https://old.reddit.com/r/Jokes/comments/4pp3no/where_did_abraham_lincoln_go_in_1865/,self.jokes,,All over the wall,Where did Abraham Lincoln go in 1865?,2
post,4pp2th,2qh72,jokes,false,1466800600,https://old.reddit.com/r/Jokes/comments/4pp2th/i_have_a_joke_to_tell/,self.jokes,,Can you reddit?,I have a joke to tell.,0
post,4pp1z3,2qh72,jokes,false,1466800322,https://old.reddit.com/r/Jokes/comments/4pp1z3/the_perfect_son_a_i_have_the_perfect_son_b_does/,self.jokes,,[deleted],"The Perfect Son. A: I have the perfect son. B: Does he smoke? A: No, he doesn't. B: Does he drink whiskey? A: No, he doesn't. B: Does he ever come home late? A: No, he doesn't. B: I guess you really do have the perfect son. How old is he? A: He will be six months old next Wednesday.",1
post,4pp1yc,2qh72,jokes,false,1466800314,https://old.reddit.com/r/Jokes/comments/4pp1yc/a_bear_was_in_the_forest/,self.jokes,,"taking a dump when a rabbit walked by. The bear said, ""Hey rabbit, does shit stick to your fur?""

""No,"" replied the rabbit.

The bear picked up the rabbit and wiped his ass with him.",A bear was in the forest,6
post,4pp1nw,2qh72,jokes,false,1466800220,https://old.reddit.com/r/Jokes/comments/4pp1nw/what_jokes_doesntdont_make_any_sense_of_theyre/,self.jokes,,[deleted],What Joke(s) doesn't/don't make any sense of they're translated to english.,1
post,4pp12r,2qh72,jokes,false,1466800028,https://old.reddit.com/r/Jokes/comments/4pp12r/im_in_sticker/,self.jokes,,"I walked around with an ""I'm Out"" sticker yesterday and expected dirty looks, instead a few men winked at me and one even grabbed my bum. ","""I'm in"" sticker...",2
post,4pp0wf,2qh72,jokes,false,1466799970,https://old.reddit.com/r/Jokes/comments/4pp0wf/the_pound_is_weaker/,self.jokes,,Does that mean I lost weight?,The pound is weaker,1
post,4pp0w1,2qh72,jokes,false,1466799966,https://old.reddit.com/r/Jokes/comments/4pp0w1/q_why_doesnt_japan_have_feminists/,self.jokes,,A: Because they still hunt whales over there.,Q: Why doesn't Japan have feminists?,1
post,4pp0lu,2qh72,jokes,false,1466799869,https://old.reddit.com/r/Jokes/comments/4pp0lu/how_do_you_make_a_shortcut/,self.jokes,,With small scissors.,How do you make a shortcut?,28
post,4pp0kz,2qh72,jokes,false,1466799857,https://old.reddit.com/r/Jokes/comments/4pp0kz/rpolitics/,self.jokes,,[removed],/r/politics,1
post,4pp0ka,2qh72,jokes,false,1466799851,https://old.reddit.com/r/Jokes/comments/4pp0ka/whats_an_even_better_way_of_losing_pounds_than/,self.jokes,,[deleted],What's an even better way of losing pounds than P90X?,0
post,4pozl4,2qh72,jokes,false,1466799516,https://old.reddit.com/r/Jokes/comments/4pozl4/a_man_sits_quietly_at_a_bar_having_a_beer/,self.jokes,,"... When the doors to the bar fly open and an old, dirty, scraggly bearded man walks in. He looks around the bar until he spots the man at the bar, quietly drinking a beer.

""You!"" The old man points at the man at the bar, ""I fucked your mother!""

The whole bar takes notice, and looks at the young man, who is still sitting at the bar quietly enjoying a beer. 

The old man takes two steps closer, points out the man at the bar again ""YOOOOOU! Your mom sucked my cock!""

Now, everyone in the bar is getting excited to possibly see a fight. They look at the man at the bar, and he is still quietly enjoying his beer. 

The old man moves even closer, pushes the younger man in the back and says ""YOOOOOOOOOU!!""

The man at the bar interrupts him, ""Dad, you're drunk. Go home.""","A man sits quietly at a bar, having a beer...",38
post,4pozat,2qh72,jokes,false,1466799417,https://old.reddit.com/r/Jokes/comments/4pozat/best_eu_jokes/,self.jokes,,[deleted],Best EU jokes?,2
post,4poz7b,2qh72,jokes,false,1466799386,https://old.reddit.com/r/Jokes/comments/4poz7b/a_scotsman_a_briton_and_claudia_schiffer_on_a/,self.jokes,,[deleted],"A Scotsman, a Briton, and Claudia Schiffer on a train...",3
post,4poysx,2qh72,jokes,false,1466799252,https://old.reddit.com/r/Jokes/comments/4poysx/what_does_the_maffia_and/,self.jokes,,"...eating pussy have in common?    
                                                               
One slip of the tongue and you're in deep shit.",What does the Maffia and...,3
post,4poyfs,2qh72,jokes,false,1466799118,https://old.reddit.com/r/Jokes/comments/4poyfs/the_british_pound_is_losing_value_so_fast/,self.jokes,,...so fast that they're renaming it the tonne to give the impression it still has weight.,The British pound is losing value so fast...,1
post,4poyd8,2qh72,jokes,false,1466799093,https://old.reddit.com/r/Jokes/comments/4poyd8/if_i_had_a_pound_for_every_brexit_joke_on_here/,self.jokes,,I'd still only have about 5 cents.,If i had a pound for every 'Brexit' joke on here...,99
post,4poxww,2qh72,jokes,false,1466798946,https://old.reddit.com/r/Jokes/comments/4poxww/a_milkman_heads_to_a_nearby_school_after_an/,self.jokes,,His milkshake really did bring the boys to the yard.,A Milkman heads to a nearby school after an Earthquake...,0
post,4poxaz,2qh72,jokes,false,1466798744,https://old.reddit.com/r/Jokes/comments/4poxaz/what_do_you_call_the_british_currency_now/,self.jokes,,[deleted],What do you call the British currency now?,0
post,4poxar,2qh72,jokes,false,1466798743,https://old.reddit.com/r/Jokes/comments/4poxar/what_do_you_get_if_you_insert_human_dna_into_a/,self.jokes,,[deleted],What do you get if you insert human DNA into a goat?,56
post,4powxb,2qh72,jokes,false,1466798626,https://old.reddit.com/r/Jokes/comments/4powxb/why_cant_you_hear_a_pterodactyl_using_the_restroom/,self.jokes,,Because they're extinct ,Why can't you hear a pterodactyl using the restroom?,75
post,4powhb,2qh72,jokes,false,1466798480,https://old.reddit.com/r/Jokes/comments/4powhb/donald_trump_hillary_clinton_and_a_voter_walk/,self.jokes,,[deleted],"Donald Trump, Hillary Clinton, and a Voter walk into a bar...",6
post,4pow8o,2qh72,jokes,false,1466798394,https://old.reddit.com/r/Jokes/comments/4pow8o/three_british_nuns_die_in_a_car_crash/,self.jokes,,"They arrive to The Gates, where St Peter awaits for them:

""Ah, you've arrived my daughters! Please have no fear, for you are nuns and will surely go to heaven. But before that, you must confess your sins and wash any sin off your body.""

They form a queue and the first takes a step forward and says,

- I confess! I have, once in a lifetime, masturbated a man!

- Well then, says Peter, wash your hands in this holy basin of water.

As she does so, an argument breaks out between the other two. Intrigued, Peter asks what the problem is.

I would like to wash my mouth before the other one washes her buttocks, says the last in line.

edit: grammar ",Three British Nuns Die in a Car Crash,0
post,4poucp,2qh72,jokes,false,1466797749,https://old.reddit.com/r/Jokes/comments/4poucp/what_did_the_prostitute_wear_under_her_bikini/,self.jokes,,[deleted],What did the prostitute wear under her bikini bottom?,1
post,4pou2e,2qh72,jokes,false,1466797657,https://old.reddit.com/r/Jokes/comments/4pou2e/what_did_the_sheep_say_to_the_farmers_crop/,self.jokes,,This is baaaad. ,What did the sheep say to the farmers crop?,1
post,4pot5v,2qh72,jokes,false,1466797363,https://old.reddit.com/r/Jokes/comments/4pot5v/i_dont_understand_why_people_are_so_amazed_when_i/,self.jokes,,[removed],"I don't understand why people are so amazed when I say my grandfather survived Auschwitz. I mean, most German Officers did.",1
post,4posvt,2qh72,jokes,false,1466797279,https://old.reddit.com/r/Jokes/comments/4posvt/a_kid_woks_up_to_his_teachir_with_a_nife/,self.jokes,,[removed],A kid woks up to his teachir with a nife!,1
post,4poskp,2qh72,jokes,false,1466797177,https://old.reddit.com/r/Jokes/comments/4poskp/a_police_officer_on_a_bike_route_sees_2_men/,self.jokes,,"The officer slows down to observe, and to see if the argument would become violent. The 2 men are bitter, and get louder by the minute. Suddenly, they both reach into their pockets. The first man pulls out some sodium chloride and throws it at the second man, while the second man get a 9 volt and 2 AA's and throws them at the first man.

The officer calls for backup, and the 2 men are arrested for assault and battery.",A police officer on a bike route sees 2 men arguing.,5
post,4poshu,2qh72,jokes,false,1466797152,https://old.reddit.com/r/Jokes/comments/4poshu/british_food_and_british_women/,self.jokes,,[deleted],British food and British women,0
post,4pos1f,2qh72,jokes,false,1466797009,https://old.reddit.com/r/Jokes/comments/4pos1f/i_just_found_out_diarrhea_is_genetic/,self.jokes,,It runs in your genes.,I just found out diarrhea is genetic...,24
post,4porv3,2qh72,jokes,false,1466796950,https://old.reddit.com/r/Jokes/comments/4porv3/today_i_got_my_first_period/,self.jokes,,pay period. CHOOM!,Today I got my first period...,0
post,4pornb,2qh72,jokes,false,1466796882,https://old.reddit.com/r/Jokes/comments/4pornb/an_airplane_carrying_pepsi_crashes/,self.jokes,,"An airplane full of a shipment of Pepsi flying over Africa had a malfunction, and went down. A few weeks later, the Pepsi Company sent a rescue plane. They searched the area and found a tribe of cannibals. 

They walked up to the Chief of the tribe and asked him if he knew anything about the crash. 

The Chief said, ""You betcha!"" 

When asked where the crew was, the Chief replied, ""We ate the crew, and we drank the Pepsi."" 

The Rescue crew were shocked. One man asked, ""Did you eat their legs?"" 

The chief replied, ""We ate their legs, and we drank the Pepsi."" 

Another rescuer asked, ""Did you eat their arms?"" 

The Chief replied, ""We ate their arms, and we drank the Pepsi."" 

After looking totally perplexed for a minute, a third asked, ""Did you...you know...eat, their...'things'?"" 

The chief says, ""No."" 

""No?"" asked the rescuer. 

""No,"" replied the Chief, ""THINGS go better with Coke.""",An Airplane Carrying Pepsi Crashes...,7
post,4porl2,2qh72,jokes,false,1466796865,https://old.reddit.com/r/Jokes/comments/4porl2/just_got_my_first_ever_gig_its_gonna_be_in_a/,self.jokes,,"Im playing the triangle, me stand at the back an ting","Just got my first ever gig, its gonna be in a reggae band.",0
post,4poqym,2qh72,jokes,false,1466796665,https://old.reddit.com/r/Jokes/comments/4poqym/i_was_stood_in_line_at_tescos_earlier_today/,self.jokes,,"...and there was a foreign couple in front of me checking out. The cashier asked them if they'd like any help packing their bags, and I thought 'blimey, that's happening quickly!'",I was stood in line at Tesco's earlier today...,1
post,4poqp4,2qh72,jokes,false,1466796590,https://old.reddit.com/r/Jokes/comments/4poqp4/the_united_kingdom/,self.jokes,,[removed],The United Kingdom,1
post,4poqjn,2qh72,jokes,false,1466796537,https://old.reddit.com/r/Jokes/comments/4poqjn/steve_martin_green_lights_female_cast_remake_of/,self.jokes,,Apparently my wife got the lead role.,"Steve Martin green lights female cast remake of ""The Jerk"" called ""The Bitch""",0
post,4poqb4,2qh72,jokes,false,1466796457,https://old.reddit.com/r/Jokes/comments/4poqb4/sitting_on_the_toilet/,self.jokes,,Scrolling through dating apps while on the toilet is the best idea... etiher way you're gonna find shit.,Sitting on the Toilet,3
post,4poq41,2qh72,jokes,false,1466796393,https://old.reddit.com/r/Jokes/comments/4poq41/when_do_jewish_people_believe_the_fetus_achieves/,self.jokes,,"Not until he graduates from medical school. 

Heard this one from a Jewish patient I had once. ",When do Jewish people believe the fetus achieves viability?,2
post,4popej,2qh72,jokes,false,1466796166,https://old.reddit.com/r/Jokes/comments/4popej/til_a_russian_match_official_was_once_jailed_for/,self.jokes,,oops wrong sub,TIL A Russian Match Official was once jailed for making the wrong substitution at a world cup match,0
post,4popbl,2qh72,jokes,false,1466796137,https://old.reddit.com/r/Jokes/comments/4popbl/in_a_way_im_happy_that_brexit_happened/,self.jokes,,Now I don't need to correct people when they refer to the UK as England.,"In a way, I'm happy that Brexit happened.",3
post,4pop4t,2qh72,jokes,false,1466796077,https://old.reddit.com/r/Jokes/comments/4pop4t/a_guy_goes_to_the_doctor_doc_i_cant_stop_singing/,self.jokes,,[removed],"A guy goes to the doctor. ""Doc, I can't stop singing 'Sex Bomb.'""",1
post,4pop3j,2qh72,jokes,false,1466796065,https://old.reddit.com/r/Jokes/comments/4pop3j/my_girlfriend_told_me_if_this_get_200_upvotes_we/,self.jokes,,Please don't upvote her strap on is huge!,My Girlfriend told me if this get 200 upvotes we would try anal,0
post,4poop2,2qh72,jokes,false,1466795936,https://old.reddit.com/r/Jokes/comments/4poop2/steve_martin_green_lights_female_cast_remake_of/,self.jokes,,[deleted],"Steve Martin green lights female cast remake of ""The Jerk"" called ""The Bitch""",1
post,4poolt,2qh72,jokes,false,1466795907,https://old.reddit.com/r/Jokes/comments/4poolt/what_do_you_get_when_you_piss_off_the_avengers/,self.jokes,,Nick's fury.,What do you get when you piss off the Avengers?,0
post,4poo2m,2qh72,jokes,false,1466795741,https://old.reddit.com/r/Jokes/comments/4poo2m/im_training_for_a_marathon_with_my_friend_every/,self.jokes,,It's a running joke.,"I'm training for a marathon with my friend. Every day when we hit the trails he tells me the same thing, and it always makes me laugh.",16
post,4ponrz,2qh72,jokes,false,1466795639,https://old.reddit.com/r/Jokes/comments/4ponrz/did_you_hear_about_the_new_brexit_diet/,self.jokes,,You do something incredibly stupid and you lose pounds fast.,Did you hear about the new Brexit diet?,0
post,4pongr,2qh72,jokes,false,1466795546,https://old.reddit.com/r/Jokes/comments/4pongr/do_i_look_thinner_to_you/,self.jokes,,[deleted],Do I look thinner to you?,1
post,4ponec,2qh72,jokes,false,1466795522,https://old.reddit.com/r/Jokes/comments/4ponec/too_long_a_title_joke_is_below/,self.jokes,,[removed],"Too long a title, joke is below:",1
post,4pomfc,2qh72,jokes,false,1466795212,https://old.reddit.com/r/Jokes/comments/4pomfc/i_like_my_stock_market_the_way_i_like_my_airplanes/,self.jokes,,[deleted],I like my Stock Market the way I like my Airplanes,0
post,4pomaj,2qh72,jokes,false,1466795169,https://old.reddit.com/r/Jokes/comments/4pomaj/whole_joke_inside/,self.jokes,,"An arab walks in to a gay bar. The bar tender asks ""What are you havin?""

""Shots for everyone!""",whole joke inside,0
post,4polyf,2qh72,jokes,false,1466795069,https://old.reddit.com/r/Jokes/comments/4polyf/a_funny_joke_is_below_this_sentence/,self.jokes,,"                                        
                                This sentence
                       _______________________
                                  A funny joke
",A funny joke is below this sentence.,0
post,4polw3,2qh72,jokes,false,1466795053,https://old.reddit.com/r/Jokes/comments/4polw3/what_word_that_starts_with_an_n_and_ends_with_an/,self.jokes,,Neighbor,"What word that starts with an ""N"" and ends with an ""R"" would you never want to call a black person",27
post,4polqk,2qh72,jokes,false,1466795006,https://old.reddit.com/r/Jokes/comments/4polqk/dad_can_i_borrow_10_pounds/,self.jokes,,- 15 pounds? Why do you need 20 pounds?,"- Dad, can I borrow 10 pounds?",404
post,4polnu,2qh72,jokes,false,1466794985,https://old.reddit.com/r/Jokes/comments/4polnu/britain_best_strike_a_deal_with_magic_stars_dont/,self.jokes,,"Yes

",Britain best strike a deal with magic stars. don't screw me twice in one day world.,0
post,4pol4t,2qh72,jokes,false,1466794831,https://old.reddit.com/r/Jokes/comments/4pol4t/one_could_say_that_brexit_has_been/,self.jokes,,... quite secessful.,One could say that Brexit has been ...,15
post,4pol2j,2qh72,jokes,false,1466794809,https://old.reddit.com/r/Jokes/comments/4pol2j/whats_the_name_of_the_national_ethipian_sea_animal/,self.jokes,,A starvefish,What's the name of the national Ethipian sea animal?,0
post,4poktl,2qh72,jokes,false,1466794727,https://old.reddit.com/r/Jokes/comments/4poktl/what_do_you_call_a_three_humped_camel/,self.jokes,,"I don't ... know ... what?

Pregnant.

hahahaha.",What do you call a three humped camel?,0
post,4pokq5,2qh72,jokes,false,1466794702,https://old.reddit.com/r/Jokes/comments/4pokq5/wanna_hear_a_joke/,self.jokes,,[deleted],Wanna hear a joke?,2
post,4pokdc,2qh72,jokes,false,1466794572,https://old.reddit.com/r/Jokes/comments/4pokdc/brexit/,self.jokes,,[removed],Brexit.,1
post,4pojek,2qh72,jokes,false,1466794245,https://old.reddit.com/r/Jokes/comments/4pojek/how_babies_are_made/,self.jokes,,[deleted],How babies are made?,0
post,4poj8o,2qh72,jokes,false,1466794200,https://old.reddit.com/r/Jokes/comments/4poj8o/islam_is_a_religion_of_peace/,self.jokes,,[removed],Islam is a religion of peace.,1
post,4poikm,2qh72,jokes,false,1466793993,https://old.reddit.com/r/Jokes/comments/4poikm/the_uks_referendum_on_eu_membership_sponsored_by/,self.jokes,,What's the worst that could happen? ,"The UK's referendum on EU membership, sponsored by Dr. Pepper",0
post,4poi7d,2qh72,jokes,false,1466793874,https://old.reddit.com/r/Jokes/comments/4poi7d/great_britain_voted_brexit/,self.jokes,,[deleted],Great Britain voted Brexit...,0
post,4pohtw,2qh72,jokes,false,1466793753,https://old.reddit.com/r/Jokes/comments/4pohtw/earlier_today_in_a_supermarket_in_the_uk_the/,self.jokes,,"Earlier today in a supermarket in the UK, the cashier asked the Foreign couple in front of me if they wanted help packing their bags. Fuck me, we only voted out yesterday, give them a chance!",Earlier today in a supermarket in the UK the cashier asked the...,1
post,4pohmk,2qh72,jokes,false,1466793687,https://old.reddit.com/r/Jokes/comments/4pohmk/where_do_german_parents_send_their_add_kids/,self.jokes,,Concentration Camps,Where do german parents send their ADD kids?,271
post,4pohh0,2qh72,jokes,false,1466793633,https://old.reddit.com/r/Jokes/comments/4pohh0/murica/,self.jokes,,[deleted],Murica...,1
post,4poh0y,2qh72,jokes,false,1466793496,https://old.reddit.com/r/Jokes/comments/4poh0y/wanna_hear_a_joke/,self.jokes,,[deleted],Wanna hear a joke?,1
post,4pogwt,2qh72,jokes,false,1466793458,https://old.reddit.com/r/Jokes/comments/4pogwt/brexit/,self.jokes,,[removed],Brexit,1
post,4pogj7,2qh72,jokes,false,1466793351,https://old.reddit.com/r/Jokes/comments/4pogj7/a_priest_and_a_ny_cab_driver_died_together_and/,self.jokes,,"A Priest and a NY Cab Driver died together and went to heaven. They get to the pearly gates and an angel greets them. First the angel takes them to the NY cab drivers house in heaven. It's amazing it has marble floors a butler and maid and a swimming pool it's awesome, the Cab drivers thanks the angel and they move on to the priest's residence. Needless to say it's a log cabin with no water or electricity. The priest is amazed at the simple house compared to the NY cab driver and he bursts out at the angle and says how could this be I spent my entire life dedicated to g-d. The angel responds it's simple. Every sunday you would go up and give a sermon and everyone fell asleep, but when this NY cab driver drove everyone prayed!!.",A Priest and a NY Cab Driver died together and went to heaven,25
post,4pogiy,2qh72,jokes,false,1466793349,https://old.reddit.com/r/Jokes/comments/4pogiy/what_did_mike_tyson_say_to_vincent_van_gogh/,self.jokes,,You gonna eat that?,What did Mike Tyson say to Vincent Van Gogh?,84
post,4pogdo,2qh72,jokes,false,1466793300,https://old.reddit.com/r/Jokes/comments/4pogdo/why_does_the_chicken_coop_have_2_doors/,self.jokes,,[deleted],Why does the chicken coop have 2 doors?,0
post,4pogdb,2qh72,jokes,false,1466793298,https://old.reddit.com/r/Jokes/comments/4pogdb/how_do_we_know_that_adam_wasnt_a_black_man/,self.jokes,,Have you ever tried taking a rib from a black man!!?!,How do we know that Adam wasn't a black man?,12
post,4pog3j,2qh72,jokes,false,1466793224,https://old.reddit.com/r/Jokes/comments/4pog3j/little_johnny_and_god/,self.jokes,,[deleted],Little Johnny and God,5
post,4pofz9,2qh72,jokes,false,1466793189,https://old.reddit.com/r/Jokes/comments/4pofz9/whats_the_difference_between_a_sociopath_and_a/,self.jokes,,[deleted],What's the difference between a sociopath and a psychopath?,1
post,4pofxb,2qh72,jokes,false,1466793168,https://old.reddit.com/r/Jokes/comments/4pofxb/im_a_cock_slut/,self.jokes,,[deleted],Im a cock slut,0
post,4pof05,2qh72,jokes,false,1466792880,https://old.reddit.com/r/Jokes/comments/4pof05/a_man_has_a_conversation_with_god/,self.jokes,,"Man: How much is a minute to you?

God: A thousand years

Man: Wow really? Ok then how much is 10 million dollars to you?

God: A penny

Man: Wow that's amazing, is it ok if I can have one of your pennies?

God: Sure thing, just give me a minute
",A man has a conversation with God,40
post,4poey0,2qh72,jokes,false,1466792860,https://old.reddit.com/r/Jokes/comments/4poey0/why_do_white_people_like_mayo/,self.jokes,,They can relate to it,Why do white people like mayo?,0
post,4poeod,2qh72,jokes,false,1466792772,https://old.reddit.com/r/Jokes/comments/4poeod/i_was_at_morrisons_earlier_and_the_cashier_asked/,self.jokes,,"I thought ""Fuck me, this is getting serious""",I was at Morrisons earlier and the cashier asked a foreign couple if they needed help packing.,6
post,4poek7,2qh72,jokes,false,1466792735,https://old.reddit.com/r/Jokes/comments/4poek7/i_like_my_women_how_i_like_my_steak/,self.jokes,,[deleted],I like my women how I like my steak.,5
post,4poefb,2qh72,jokes,false,1466792699,https://old.reddit.com/r/Jokes/comments/4poefb/what_is_the_best_thing_about_switzerland/,self.jokes,,[removed],What is the best thing about Switzerland?,1
post,4poeb2,2qh72,jokes,false,1466792663,https://old.reddit.com/r/Jokes/comments/4poeb2/whats_mr_ts_favorite_holiday/,self.jokes,,"April, Fools. ",What's Mr. T's favorite holiday?,8
post,4poe8z,2qh72,jokes,false,1466792640,https://old.reddit.com/r/Jokes/comments/4poe8z/if_you_are_moving_a_piano_from_high_storage_and/,self.jokes,,[removed],"If you are moving a piano from high storage and have the choice of using a ladder or a forklift, I would recommend the latter.",1
post,4podw3,2qh72,jokes,false,1466792524,https://old.reddit.com/r/Jokes/comments/4podw3/which_american_state_is_not_great_but_not_bad/,self.jokes,,OK.,"Which American state is not great, but not bad either?",102
post,4podsl,2qh72,jokes,false,1466792496,https://old.reddit.com/r/Jokes/comments/4podsl/a_man_comes_home_to_his_wife/,self.jokes,,"""honey,"" he says, ""pack your bags. I just won the lottery!""

""That's amazing! What should I pack?""

""I don't care. Just pack your bags and get the fuck out of here.""",A man comes home to his wife,21
post,4podet,2qh72,jokes,false,1466792396,https://old.reddit.com/r/Jokes/comments/4podet/im_addicted_to_drinking_brake_fluid/,self.jokes,,"But, I can stop whenever I want.",I'm addicted to drinking brake fluid.,511
post,4poddz,2qh72,jokes,false,1466792389,https://old.reddit.com/r/Jokes/comments/4poddz/what_is_a_pirates_favorite_subreddit_to_subscribe/,self.jokes,,[removed],What is a pirate's favorite Subreddit to subscribe to?,1
post,4pocxc,2qh72,jokes,false,1466792257,https://old.reddit.com/r/Jokes/comments/4pocxc/the_british_pound_has_lose_to_much_of_its_worth/,self.jokes,,"it will have to be renamed, the Ounce.",The British Pound has lose to much of its worth in the market crash,0
post,4pocuh,2qh72,jokes,false,1466792240,https://old.reddit.com/r/Jokes/comments/4pocuh/what_does_it_take_to_impregnate_mother_russia/,self.jokes,,[deleted],What does it take to impregnate Mother Russia?,4
post,4pocrf,2qh72,jokes,false,1466792215,https://old.reddit.com/r/Jokes/comments/4pocrf/so_i_saw_this_bear_doing_a_downward_dog_the_other/,self.jokes,,Guess you can call him Yogi Bear. ,So I saw this bear doing a downward dog the other day.,0
post,4pochl,2qh72,jokes,false,1466792124,https://old.reddit.com/r/Jokes/comments/4pochl/how_do_you_turn_an_unsubsidized_loan_into_a/,self.jokes,,Grow corn (ethanol) on it.,How do you turn an unsubsidized loan into a subsidized loan?,0
post,4poce4,2qh72,jokes,false,1466792093,https://old.reddit.com/r/Jokes/comments/4poce4/with_the_way_britain_is_going/,self.jokes,,The pound is looking more like the ounce.,With the way Britain is going...,0
post,4pocdj,2qh72,jokes,false,1466792089,https://old.reddit.com/r/Jokes/comments/4pocdj/what_is_the_difference_between_a_snowman_and_a/,self.jokes,,Snowballs.,What is the difference between a snowman and a snowwoman?,1
post,4pobv3,2qh72,jokes,false,1466791920,https://old.reddit.com/r/Jokes/comments/4pobv3/a_study_of_married_women_showed_that_90_of/,self.jokes,,The other 10% have dumb wives.,A study of married women showed that 90% of married men still masturbate,35
post,4poaiv,2qh72,jokes,false,1466791518,https://old.reddit.com/r/Jokes/comments/4poaiv/webmd_gave_me_cancer/,self.jokes,,"One don't simply leave Web Md, without getting a cancer !",WebMd. gave me Cancer !!,0
post,4poa5c,2qh72,jokes,false,1466791412,https://old.reddit.com/r/Jokes/comments/4poa5c/what_do_you_call_popcorn_laying_on_the_floor/,self.jokes,,[deleted],What do you call popcorn laying on the floor?,0
post,4po9k9,2qh72,jokes,false,1466791243,https://old.reddit.com/r/Jokes/comments/4po9k9/i_dont_know_why_everyone_is_freaking_out_about/,self.jokes,,[deleted],I don't know why everyone is freaking out about the Brexit.,1
post,4po99m,2qh72,jokes,false,1466791157,https://old.reddit.com/r/Jokes/comments/4po99m/whats_globally_powerful_traditionally_had_a_white/,self.jokes,,[deleted],"What's globally powerful, traditionally had a white population, but became significantly more diverse after losing 1GB?",0
post,4po984,2qh72,jokes,false,1466791142,https://old.reddit.com/r/Jokes/comments/4po984/a_man_walked_up_to_me_on_the_street_and_handed_me/,self.jokes,,I couldn't believe he was able to check my battery so quickly...,"A man walked up to me on the street and handed me a flyer that said ""Free car-battery check, no charge.""",3
post,4po8yl,2qh72,jokes,false,1466791062,https://old.reddit.com/r/Jokes/comments/4po8yl/britain_should_have_written_a_break_up_note/,self.jokes,,"""It's not EU, it's me""",Britain should have written a break up note,262
post,4po8t2,2qh72,jokes,false,1466791010,https://old.reddit.com/r/Jokes/comments/4po8t2/2016/,self.jokes,,[removed],2016,1
post,4po8ek,2qh72,jokes,false,1466790879,https://old.reddit.com/r/Jokes/comments/4po8ek/what_do_you_call_a_friendly_helicopter/,self.jokes,,A hello-copter,What do you call a friendly helicopter?,3
post,4po81p,2qh72,jokes,false,1466790760,https://old.reddit.com/r/Jokes/comments/4po81p/what_do_you_tell_a_woman_with_two_black_eyes/,self.jokes,,Nothing! You already told her twice!!,What do you tell a woman with two black eyes?,0
post,4po80l,2qh72,jokes,false,1466790752,https://old.reddit.com/r/Jokes/comments/4po80l/i_had_a_dream_last_night/,self.jokes,,That a hamburger was eating  me!,I had a dream last night...,0
post,4po800,2qh72,jokes,false,1466790747,https://old.reddit.com/r/Jokes/comments/4po800/what_do_pubes_and_salad_have_in_common/,self.jokes,,[deleted],What do pubes and salad have in common?,12
post,4po7yd,2qh72,jokes,false,1466790731,https://old.reddit.com/r/Jokes/comments/4po7yd/i_stopped_a_kidnapping_today/,self.jokes,,I woke him up,I stopped a kidnapping today..,25
post,4po7a0,2qh72,jokes,false,1466790516,https://old.reddit.com/r/Jokes/comments/4po7a0/wasnt_by_british_accent_great/,self.jokes,,I thought all British accents were Great British accents,Wasn't by British accent great?,0
post,4po76v,2qh72,jokes,false,1466790488,https://old.reddit.com/r/Jokes/comments/4po76v/what_will_be_the_name_of_a_movie_where_all/,self.jokes,,No country for old woman.,What will be the name of a movie where all countries of UK decides to leave UK?,0
post,4po74f,2qh72,jokes,false,1466790470,https://old.reddit.com/r/Jokes/comments/4po74f/what_separates_man_from_animals/,self.jokes,,"According to Donald Trump, the wall he is going to build.",What separates man from animals?,18
post,4po6bq,2qh72,jokes,false,1466790222,https://old.reddit.com/r/Jokes/comments/4po6bq/a_jewish_man_trying_to_win_the_lottery/,self.jokes,,"A Jewish man in Israel goes to the Western Wall every day for 25 years and puts a note saying ""Please let me win the lottery"". One day he goes, God is looking down at him post the note. ""God, he's been coming here for 25 years posting the same note and hasn't missed a day. Why not let him win the lottery?"" says God's assistant. God says ""I will, once he actually starts playing"".",A Jewish man trying to win the lottery.,0
post,4po68s,2qh72,jokes,false,1466790194,https://old.reddit.com/r/Jokes/comments/4po68s/claustrophobic_people_are_interesting/,self.jokes,,Because they always try to think outside of the box.,Claustrophobic people are interesting,9
post,4po65t,2qh72,jokes,false,1466790167,https://old.reddit.com/r/Jokes/comments/4po65t/how_do_you_torture_a_british_person/,self.jokes,,[deleted],how do you torture a british person?,0
post,4po63p,2qh72,jokes,false,1466790148,https://old.reddit.com/r/Jokes/comments/4po63p/i_have_a_lumberjack_funny_for_yall/,self.jokes,,"One lumberjack asks ""why are we cutting down all these trees?"" The other one says ""for profit, AND competition"". The first lumberjack asks, ""but isn't that wrong, and detrimental to the environment?"" And then they chopped all the trees down and we all suffocated BECAUSE without trees, humans would not be able survive because the air would be bad for breathing. If anything, people would have to develop gas masks that filter the little oxygen that would be left in the air. Trees are a crucial part of the carbon cycle, a global process in which carbon dioxide constantly circulates through the atmosphere into organism and back again LOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOLOL!!!!",I have a Lumberjack funny for yall.,0
post,4po61i,2qh72,jokes,false,1466790131,https://old.reddit.com/r/Jokes/comments/4po61i/i_walked_into_a_gay_bar_full_of_colorful_gay_men/,self.jokes,,[deleted],I walked into a gay bar full of colorful gay men masturbating,0
post,4po5um,2qh72,jokes,false,1466790074,https://old.reddit.com/r/Jokes/comments/4po5um/so_there_was_a_guy_who/,self.jokes,,",after a long day of driving, wanted to find a  place to sleep. After driving for a while he came across a small farm. Thinking oh well it can't be that bad he knocks on the door and asks the man if he can spend the night at his farm. The man says yes on one condition ""you cannot go into my cellur"". The man just wanting to sleeps accepts this condition and goes to his room. Later that night the man can't sleep because he can't stop thinking about what in the world could be down in his cellur. After hours of thinking he finally gets up from his bed and goes to investigate. He goes down into the cellur and in the center is a cage with a purple gorilla in it and a sign next to it saying do not touch. Hmm well already breaking the other rule the man decides he wants to know what a purple gorilla would feel like. So he reaches in and touches it. As soon as he does the gorilla goes ape shit crazy. It begins yelling and screaming trying to reach out for the man through the bars. Unable to reach him  the gorilla grabs the bars and using an immense amout of strength bends them open. The man, scared out of goddamn mind,immedietly runs up stairs and gets in his truck and begins driving. He starts going 40 miles an hour and bam there was the gorilla right behind so he starts to speed up to 60 70 80 miles per hour and to no avail the gorilla is still hot on his tail. Suddenly the gorilla jumps up onto the back of the truck. He grabs the windows and tears them off with an ungodly amount of strength. Suddenly the gorilla reaches through and touches the man's shoulder and says ""Your it"".",So there was a guy who,2
post,4po59j,2qh72,jokes,false,1466789892,https://old.reddit.com/r/Jokes/comments/4po59j/remember_when_the_uk_was_part_of_the_eu/,self.jokes,,It seems like only yesterday.,Remember When the UK Was Part of the EU?,1
post,4po4r7,2qh72,jokes,false,1466789750,https://old.reddit.com/r/Jokes/comments/4po4r7/a_man_love_his_son/,self.jokes,,"a man love his son a lot but his son nothing,,,,,,,,,,",A man love his son,0
post,4po4is,2qh72,jokes,false,1466789679,https://old.reddit.com/r/Jokes/comments/4po4is/queen_reacts_to_brexit/,self.jokes,,"Bloody hell, my kingdom is in tatters! \*sips tea\*
",Queen reacts to Brexit,0
post,4po4aj,2qh72,jokes,false,1466789614,https://old.reddit.com/r/Jokes/comments/4po4aj/a_feminist_once_asked_me_how_i_viewed_lesbians/,self.jokes,,[deleted],A feminist once asked me how I viewed lesbians.,27
post,4po3m9,2qh72,jokes,false,1466789410,https://old.reddit.com/r/Jokes/comments/4po3m9/so_many_british_jokes_after_the_brexit_vote/,self.jokes,,"EU, it's disgusting.

At least I tried",So many British jokes after the Brexit Vote.,1
post,4po39m,2qh72,jokes,false,1466789293,https://old.reddit.com/r/Jokes/comments/4po39m/what_kind_of_bagel_can_fly/,self.jokes,,A plain bagel.,What kind of bagel can fly?,1
post,4po2td,2qh72,jokes,false,1466789153,https://old.reddit.com/r/Jokes/comments/4po2td/an_old_arab_in_the_usa_wants_to_plant_potatoes/,self.jokes,,"... but being the old age that he is, he cannot. He is sad, so he writes  an e-mail to his son, whose studying in London.
 ""Hello, Ahmad, I'm sad. I'd want to plant potatoes, but I'm old and weak""
The son replies soon:
""DAD, DO NOT DIG IN THE GARDEN!! YOU'LL FIND THE THING!!!""

A week passes, and FBI agents arrive at his house. They dig through every centimetre in the garden, but they found nothing. They leave. The old arab wants to write his son about what happened,when he finds an e-mail from him.

""Hello father, your garden is probably prepared for potatoes. That's all I can do from here. Bye, Ahmad.""

E: sorry for spelling, english is my 2nd language
","An old arab in the USA want's to plant potatoes,...",28
post,4po2hc,2qh72,jokes,false,1466789041,https://old.reddit.com/r/Jokes/comments/4po2hc/did_you_know_was_a_mute_nazi_running_a/,self.jokes,,[deleted],Did you know was a mute Nazi running a concentration camp during WW2?,0
post,4po2d3,2qh72,jokes,false,1466789005,https://old.reddit.com/r/Jokes/comments/4po2d3/what_do_you_call_a_school_for_whores_that_is/,self.jokes,,A destitute institute of ill repute.,What do you call a School for Whores that is unable to pay its bills?,0
post,4po1zb,2qh72,jokes,false,1466788872,https://old.reddit.com/r/Jokes/comments/4po1zb/2016_us_presidential_elections/,self.jokes,,[removed],2016 U.S. Presidential Elections...,1
post,4po1id,2qh72,jokes,false,1466788738,https://old.reddit.com/r/Jokes/comments/4po1id/neverforget/,self.jokes,,"Wife of a Brazilian goalkeeper wakes him up: ""Honey, it's already 8!""

Him: ""What! Did Germany score another one?""",#NeverForget,0
post,4po1g2,2qh72,jokes,false,1466788717,https://old.reddit.com/r/Jokes/comments/4po1g2/what_do_star_wars_and_the_uk_have_in_common/,self.jokes,,They both abandoned the EU,What do star wars and the U.K. have in common?,23
post,4po1a8,2qh72,jokes,false,1466788664,https://old.reddit.com/r/Jokes/comments/4po1a8/whats_the_quickest_way_to_lose_100_pounds/,self.jokes,,Leave the European Union. . . Beep boop bop bam Pow!,What's the quickest way to lose 100 pounds?,0
post,4po0rg,2qh72,jokes,false,1466788504,https://old.reddit.com/r/Jokes/comments/4po0rg/the_uk_is_a_lot_like_my_last_blind_date/,self.jokes,,...both said: Leave Euw.,The UK is a lot like my last blind date...,0
post,4po0qw,2qh72,jokes,false,1466788500,https://old.reddit.com/r/Jokes/comments/4po0qw/so_a_feminist_gets_asked_out_an_a_date/,self.jokes,,[removed],So a feminist gets asked out an a date...,1
post,4po0pl,2qh72,jokes,false,1466788489,https://old.reddit.com/r/Jokes/comments/4po0pl/i_heard_a_really_good_joke_about_money_today/,self.jokes,,EU probably saw it on Reddit a THOUSAND FUCKING TIMES GOD DAMMIT,I heard a really good joke about money today.,2
post,4po0es,2qh72,jokes,false,1466788385,https://old.reddit.com/r/Jokes/comments/4po0es/im_dyslexic_and_an_atheist/,self.jokes,,[removed],I'm dyslexic and an atheist,1
post,4po0a5,2qh72,jokes,false,1466788343,https://old.reddit.com/r/Jokes/comments/4po0a5/its_the_most_rapid_drop_in_the_value_of_sterling/,self.jokes,,Since Raheem joined City,It's the most rapid drop in the value of sterling,0
post,4pnzoq,2qh72,jokes,false,1466788170,https://old.reddit.com/r/Jokes/comments/4pnzoq/me_and_my_wife_are_like_catdog/,self.jokes,,Inseparable since birth.,Me and my wife are like Catdog...,0
post,4pnzhq,2qh72,jokes,false,1466788104,https://old.reddit.com/r/Jokes/comments/4pnzhq/did_you_hear_why_santa_stopped_going_down_chimneys/,self.jokes,,He was getting Claus-trophobic.,Did you hear why Santa stopped going down Chimneys?,1
post,4pnyvc,2qh72,jokes,false,1466787894,https://old.reddit.com/r/Jokes/comments/4pnyvc/whats_rickon_starks_favourite_band/,self.jokes,,One Direction ,What's Rickon Starks favourite band?,5
post,4pnyn8,2qh72,jokes,false,1466787839,https://old.reddit.com/r/Jokes/comments/4pnyn8/whats_bill_gatess_favorite_dessert/,self.jokes,,apple turnover,What's Bill Gates's favorite dessert,16
post,4pnyfv,2qh72,jokes,false,1466787780,https://old.reddit.com/r/Jokes/comments/4pnyfv/britain_lied/,self.jokes,,[removed],Britain lied...,1
post,4pnybf,2qh72,jokes,false,1466787750,https://old.reddit.com/r/Jokes/comments/4pnybf/now_i_understand_why_the_british_population_was/,self.jokes,,Brits are really good at pulling out.,Now I understand why the British population was on a steady decline these past few years...,46
post,4pnxll,2qh72,jokes,false,1466787544,https://old.reddit.com/r/Jokes/comments/4pnxll/isnt_swallowing_semen_technically_canibalism/,self.jokes,,"I don't know, I just do it for the taste...",Isn't swallowing semen technically canibalism?,1
post,4pnxli,2qh72,jokes,false,1466787544,https://old.reddit.com/r/Jokes/comments/4pnxli/what_do_you_call_a_zombie_crossing_the_street/,self.jokes,,A Jaywalker,What do you call a zombie crossing the street?,1
post,4pnxb2,2qh72,jokes,false,1466787442,https://old.reddit.com/r/Jokes/comments/4pnxb2/why_didnt_the_england_soccer_team_didnt_vote_in/,self.jokes,,[deleted],Why didn't the England soccer team didn't vote in the EU referendum?,0
post,4pnwlj,2qh72,jokes,false,1466787226,https://old.reddit.com/r/Jokes/comments/4pnwlj/knock_knock/,self.jokes,,"""Who's there?""

""It's Britain, hurry up and answer the door.""

""Britain who?""

""Fuck this, were leaving.""",Knock knock...,2
post,4pnwg2,2qh72,jokes,false,1466787183,https://old.reddit.com/r/Jokes/comments/4pnwg2/why_did_britain_manage_the_brexit/,self.jokes,,"Most of them wanted to escape the EU, and made a break for it.",Why did Britain manage the Brexit?,0
post,4pnvxs,2qh72,jokes,false,1466787038,https://old.reddit.com/r/Jokes/comments/4pnvxs/reddit_revere/,self.jokes,,"The British are leaving, the British are leaving!",Reddit Revere,0
post,4pnv88,2qh72,jokes,false,1466786823,https://old.reddit.com/r/Jokes/comments/4pnv88/i_guess_you_could_say_europe_now_has_1_gb_of_free/,self.jokes,,[removed],I guess you could say Europe now has 1 GB of free space.,1
post,4pnutt,2qh72,jokes,false,1466786690,https://old.reddit.com/r/Jokes/comments/4pnutt/3_years_ago_i_asked_the_girl_of_my_dreams_out_and/,self.jokes,,She said no both times. ,"3 years ago I asked the girl of my dreams out, and today I asked her to marry me.",0
post,4pnuo2,2qh72,jokes,false,1466786637,https://old.reddit.com/r/Jokes/comments/4pnuo2/a_blonde_her_thermos/,self.jokes,,"A blonde notices that her coworker has a thermos, so she asks him what it's for. He responds, ""It keeps hot things hot and cold things cold.""

The blonde immediately buys one for herself. The next day, she goes to work and proudly displays it.

Her coworker asks, ""What do you have in it?""

She replies, ""Soup and ice cream.""",A Blonde &amp; Her Thermos,10
post,4pnuhu,2qh72,jokes,false,1466786579,https://old.reddit.com/r/Jokes/comments/4pnuhu/did_you_hear_the_joke_about_the_model_in_the/,self.jokes,,Never mind it was pretty shitty. ,Did you hear the joke about the model in the public restroom?,2
post,4pntow,2qh72,jokes,false,1466786322,https://old.reddit.com/r/Jokes/comments/4pntow/some_good_news_for_uk/,self.jokes,,[deleted],Some good news for UK,0
post,4pntm7,2qh72,jokes,false,1466786296,https://old.reddit.com/r/Jokes/comments/4pntm7/because_brexit/,self.jokes,,"Son: Father, I need 5 Pound for tea.

Father: 10 Pound? Why do you need 20 Pound?",Because BREXIT,0
post,4pnsuo,2qh72,jokes,false,1466786065,https://old.reddit.com/r/Jokes/comments/4pnsuo/it_is_so_hot_here/,self.jokes,,[deleted],It is so hot here...,0
post,4pns1t,2qh72,jokes,false,1466785815,https://old.reddit.com/r/Jokes/comments/4pns1t/two_jews_walk_into_a_bar/,self.jokes,,Oy Oy!,Two Jews walk into a bar...,0
post,4pnrv7,2qh72,jokes,false,1466785759,https://old.reddit.com/r/Jokes/comments/4pnrv7/the_eu_now_has_1gb_of_free_space/,self.jokes,,[removed],The EU now has 1GB of free space,1
post,4pnrhw,2qh72,jokes,false,1466785651,https://old.reddit.com/r/Jokes/comments/4pnrhw/have_you_heard_of_the_brexit_exercise/,self.jokes,,[deleted],Have you heard of the Brexit exercise?,0
post,4pnrhf,2qh72,jokes,false,1466785646,https://old.reddit.com/r/Jokes/comments/4pnrhf/i_got_a_joke_for_you/,self.jokes,,[deleted],I got a joke for you,0
post,4pnr1l,2qh72,jokes,false,1466785513,https://old.reddit.com/r/Jokes/comments/4pnr1l/todays_national_report/,self.jokes,,[deleted],Today's National Report:,0
post,4pnppa,2qh72,jokes,false,1466785082,https://old.reddit.com/r/Jokes/comments/4pnppa/how_did_the_buckets_mom_know_he_was_sick/,self.jokes,,He was a little pail.,How did the bucket's mom know he was sick?,104
post,4pnotr,2qh72,jokes,false,1466784822,https://old.reddit.com/r/Jokes/comments/4pnotr/the_leave_camp_has_picked_right_where/,self.jokes,,[deleted],The Leave camp has picked right where,0
post,4pnot1,2qh72,jokes,false,1466784816,https://old.reddit.com/r/Jokes/comments/4pnot1/what_is_the_only_job_you_can_apply_for_when_youre/,self.jokes,,[deleted],What is the only job you can apply for when you're under FBI investigation?,1
post,4pnodo,2qh72,jokes,false,1466784693,https://old.reddit.com/r/Jokes/comments/4pnodo/what_do_you_call_a_spiral_penis/,self.jokes,,[deleted],What do you call a spiral penis?,6
post,4pnod9,2qh72,jokes,false,1466784691,https://old.reddit.com/r/Jokes/comments/4pnod9/the_uk_votes_on_the_possibility_of_leaving_the_eu/,self.jokes,,It goes through,The UK votes on the possibility of leaving the EU,0
post,4pno8z,2qh72,jokes,false,1466784655,https://old.reddit.com/r/Jokes/comments/4pno8z/breaking_ongoing_kidnapping_situation_in_uk/,self.jokes,,[removed],BREAKING: Ongoing kidnapping situation in UK.,1
post,4pnnw0,2qh72,jokes,false,1466784546,https://old.reddit.com/r/Jokes/comments/4pnnw0/i_like_my_eu_like_i_like_banging_my_gf/,self.jokes,,Poundead,I like my EU like I like banging my gf...,2
post,4pnmrw,2qh72,jokes,false,1466784210,https://old.reddit.com/r/Jokes/comments/4pnmrw/the_probrexitists/,self.jokes,,can go bruck themselves.,The pro-Brexitists,0
post,4pnmqh,2qh72,jokes,false,1466784196,https://old.reddit.com/r/Jokes/comments/4pnmqh/i_guess_the_eu_has_1_gb_of_free_space_now/,self.jokes,,[removed],I guess the EU has 1 GB of free space now.,1
post,4pnmaq,2qh72,jokes,false,1466784064,https://old.reddit.com/r/Jokes/comments/4pnmaq/the_british_government_is_renaming_the_pound/,self.jokes,,They figured the ounce was more appropriate.,The British government is renaming the pound,1
post,4pnlou,2qh72,jokes,false,1466783878,https://old.reddit.com/r/Jokes/comments/4pnlou/the_uks_economy/,self.jokes,,That's the joke.,The UK's economy.,4
post,4pnl24,2qh72,jokes,false,1466783671,https://old.reddit.com/r/Jokes/comments/4pnl24/how_does_a_gay_guy_remove_a_condom/,self.jokes,,He farts,How does a gay guy remove a condom?,5
post,4pnklz,2qh72,jokes,false,1466783522,https://old.reddit.com/r/Jokes/comments/4pnklz/laying_on_my_deathbed_i_saw_life_flash_before_my/,self.jokes,,And she had some great tits!,Laying on my deathbed I saw Life flash before my eyes...,1
post,4pnk27,2qh72,jokes,false,1466783353,https://old.reddit.com/r/Jokes/comments/4pnk27/a_lumber_jack_walks_into_a_gay_bar/,self.jokes,,"It is the only bar in the small town. So the Lumber Jack figured, after a long week of work, it was going to have to do.

He walks up to the bartender and asks;

""Could I get a nice hearty lagger?""

The bartender gives a little smirk and replies;

""Certainly. Bottom or top?""

Lumber jack says;

""Tap, please.""

Bartender smiles, gives a whistle, and yells;

""Jonny Logger! You're up!""

Lumber Jack looks a little worried, so the bartender reassures him;

""Don't worry, he is the best woodworker I know. And he usually does best on top. He can fell the strongest wood, and doesn't mind it getting messy or dirty.""

Lumber Jack high tails it out of there.



Edit: Accents

Top- Tap

Bottom- Bottle

Lager- Logger

Initial sentence is just filler since I came up with it on a whim.

Sorry to post a joke without a description. Thought bottom/top would be easy enough to accent into bottle/tap.",A Lumber Jack walks into a gay bar...,0
post,4pnjyf,2qh72,jokes,false,1466783323,https://old.reddit.com/r/Jokes/comments/4pnjyf/how_much_space_is_left_in_eu/,self.jokes,,1 GB,How much space is left in EU?,7
post,4pnjw0,2qh72,jokes,false,1466783301,https://old.reddit.com/r/Jokes/comments/4pnjw0/awkward/,self.jokes,,"Nigel Farage woke up this morning. ""Yay!"" he exclaimed. He turned to his wife, pecked her on the cheek and said, ""sorry, love"" as he shoved her out the door",Awkward,0
post,4pnjqm,2qh72,jokes,false,1466783260,https://old.reddit.com/r/Jokes/comments/4pnjqm/the_uks_economy/,self.jokes,,[removed],The UK's economy.,1
post,4pnj6c,2qh72,jokes,false,1466783081,https://old.reddit.com/r/Jokes/comments/4pnj6c/european_union_now_has_1_gb_of_free_space/,self.jokes,,[removed],European Union now has 1 GB of free space!,1
post,4pnj5g,2qh72,jokes,false,1466783074,https://old.reddit.com/r/Jokes/comments/4pnj5g/fast_joke/,self.jokes,,[deleted],Fast joke.,1
post,4pnj34,2qh72,jokes,false,1466783053,https://old.reddit.com/r/Jokes/comments/4pnj34/pregnant_prostitute/,self.jokes,,"Doctor asks a pregnant prostitute, ""Do you know who the father is?""   

The prostitute  replied, ""If you ate a can of beans would you know which one made you fart?"" ",Pregnant Prostitute,2
post,4pnj1s,2qh72,jokes,false,1466783040,https://old.reddit.com/r/Jokes/comments/4pnj1s/the_ira_have_been_fighting_for_irish/,self.jokes,,All they needed to do was vote for the Conservatives. ,The IRA have been fighting for Irish reunification since the 70s. . .,9
post,4pnj0k,2qh72,jokes,false,1466783027,https://old.reddit.com/r/Jokes/comments/4pnj0k/what_the_quickest_way_to_lose_100_pounds/,self.jokes,,[deleted],What the quickest way to lose 100 pounds?,0
post,4pnijn,2qh72,jokes,false,1466782866,https://old.reddit.com/r/Jokes/comments/4pnijn/if_i_had_a_dollar_for_every_time_i_beat_off/,self.jokes,,[deleted],If I had a dollar for every time I beat off,0
post,4pnidf,2qh72,jokes,false,1466782811,https://old.reddit.com/r/Jokes/comments/4pnidf/why_do_women_wear_makeup_and_perfume/,self.jokes,,[deleted],Why do women wear makeup and perfume?,0
post,4pnhxp,2qh72,jokes,false,1466782665,https://old.reddit.com/r/Jokes/comments/4pnhxp/omg_i_just_won_the_lottery/,self.jokes,,[deleted],OMG I just won the lottery!,1
post,4pngjm,2qh72,jokes,false,1466782217,https://old.reddit.com/r/Jokes/comments/4pngjm/stupid_father/,self.jokes,,"A guy goes to the supermarket and notices an attractive woman waving at him. She says hello. He’s rather taken aback because he can’t place where he knows her from. So he says, ""Do you know me?"" To which she replies, ""I think you’re the father of one of my kids."" Now his mind travels back to the only time he has ever been unfaithful to his wife and says, ""My God, are you the stripper from my bachelor party that I made love to on the pool table with all my buddies watching while your partner whipped my butt with wet celery?"" She looks into his eyes and says calmly, ""No, I’m your son’s teacher.""",Stupid Father,3
post,4pngck,2qh72,jokes,false,1466782158,https://old.reddit.com/r/Jokes/comments/4pngck/the_british_are_dropping_pounds_faster_than_a/,self.jokes,,sorry plz kill me,The British are dropping pounds faster than a Biggest Loser contestant,0
post,4pngb4,2qh72,jokes,false,1466782141,https://old.reddit.com/r/Jokes/comments/4pngb4/i_like_my_women_like_i_like_my_coffee/,self.jokes,,[deleted],I like my women like I like my coffee,1
post,4png5f,2qh72,jokes,false,1466782091,https://old.reddit.com/r/Jokes/comments/4png5f/congrats_european_union/,self.jokes,,"On losing those pounds!! 
",CONGRATS European Union...,2
post,4png36,2qh72,jokes,false,1466782075,https://old.reddit.com/r/Jokes/comments/4png36/whats_a_word_that_starts_with_u_and_ends_with_w/,self.jokes,,Cloning.,"What's a word that starts with ""u"" and ends with ""w""?",89
post,4pnfs3,2qh72,jokes,false,1466781971,https://old.reddit.com/r/Jokes/comments/4pnfs3/to_the_remain_crowd_in_britain_come_to_canada/,self.jokes,,Half of the US is moving here soon anyhow.,"To the ""Remain"" crowd in Britain... come to Canada!",29
post,4pnfi5,2qh72,jokes,false,1466781882,https://old.reddit.com/r/Jokes/comments/4pnfi5/so_i_heard_the_workers_in_the_twin_towers_tried/,self.jokes,,Asking for an Air Kraft wasn't one of their better ideas.,So I heard the workers in the Twin Towers tried to have chocolate delivered to them by drone.,0
post,4pnffz,2qh72,jokes,false,1466781862,https://old.reddit.com/r/Jokes/comments/4pnffz/people_always_keep_making_jokes_about_how_people/,self.jokes,,He fell off of a guard tower and broke his neck.,"People always keep making jokes about how people died in the Holocaust, my grandpa died during the Holocaust.",4
post,4pnesd,2qh72,jokes,false,1466781650,https://old.reddit.com/r/Jokes/comments/4pnesd/the_eu_must_be_jewish/,self.jokes,,because it just had a brit milah.,The EU must be Jewish,0
post,4pnec8,2qh72,jokes,false,1466781510,https://old.reddit.com/r/Jokes/comments/4pnec8/my_friend_told_me_that_recycling_is_good_for_the/,self.jokes,,[deleted],My friend told me that recycling is good for the environment.,143
post,4pnebe,2qh72,jokes,false,1466781502,https://old.reddit.com/r/Jokes/comments/4pnebe/look_on_the_bright_side/,self.jokes,,The EU now has 1 GB of free space,Look on the bright side...,0
post,4pneaw,2qh72,jokes,false,1466781497,https://old.reddit.com/r/Jokes/comments/4pneaw/lets_be_respectful_of_each_others_beliefs/,self.jokes,,[deleted],Lets be respectful of each others beliefs...,0
post,4pne1d,2qh72,jokes,false,1466781409,https://old.reddit.com/r/Jokes/comments/4pne1d/the_pound/,self.jokes,,[removed],The Pound,1
post,4pndx4,2qh72,jokes,false,1466781368,https://old.reddit.com/r/Jokes/comments/4pndx4/my_current_best_joke/,self.jokes,,[deleted],My current best joke.,1
post,4pndmp,2qh72,jokes,false,1466781274,https://old.reddit.com/r/Jokes/comments/4pndmp/when_is_a_booger_not_a_booger/,self.jokes,,When it's snot.,When is a booger not a booger?,0
post,4pndlj,2qh72,jokes,false,1466781258,https://old.reddit.com/r/Jokes/comments/4pndlj/a_neutron_walks_into_a_bar/,self.jokes,,"...says, ""I'll have a pint of your best bitter please barkeep,  and your  finest scotch for a chaser."" The barman pours him his drinks, places them on the bar in front of him, and walks away. ""Just a moment my good man!"" exclaims the proton, ""You haven't charged me for my drinks! What do I owe you?""

""For you sir,"" replied the barman, ""no charge.""",A neutron walks into a bar...,2
post,4pndkx,2qh72,jokes,false,1466781252,https://old.reddit.com/r/Jokes/comments/4pndkx/how_do_you_destroy_an_empire/,self.jokes,,Brexit.,How do you destroy an empire?,0
post,4pncu9,2qh72,jokes,false,1466781009,https://old.reddit.com/r/Jokes/comments/4pncu9/looks_like_the_eu_now/,self.jokes,,[deleted],Looks like the EU now..,1
post,4pncol,2qh72,jokes,false,1466780957,https://old.reddit.com/r/Jokes/comments/4pncol/a_young_boy_had_just_gotten_his_driving_permit/,self.jokes,,"... and he asked his father, who was a minister, if they could start driving dad's car.

His father replied, ""We'll make a deal. You bring your grades up, study the Bible and get your hair cut.  Then we'll talk about it.""

After a month the boy came back and again asked his dad if he could use the car.

 The father said, ""Son, I've been real proud of you. You have brought your grades up, you've studied your bible very well. But you didn't get your hair cut!""  

The young man waited a moment and replied, ""You know dad, Samson had long hair, Moses had long hair, Noah and even Jesus had long hair...""

To which his father replied, ""Yeah, and all of them walked everywhere, on foot! ""

",A young boy had just gotten his driving permit...,46
post,4pncgw,2qh72,jokes,false,1466780888,https://old.reddit.com/r/Jokes/comments/4pncgw/what_happens_when_a_british_guy_makes_a_promise/,self.jokes,,He Brexit,What happens when a British guy makes a promise?,192
post,4pnceu,2qh72,jokes,false,1466780873,https://old.reddit.com/r/Jokes/comments/4pnceu/im_laying_in_bed_reading_a_book_when_my_dad_walks/,self.jokes,,"About five feet away from me he stops and starts pushing the tape out to me. 

It gets closer and closer until it eventually pushes against my cheek.

I ask him ""What are you doing?""

""I'm measuring your patience.""","I'm laying in bed reading a book, when my dad walks in with a tape measure...",320
post,4pnc9a,2qh72,jokes,false,1466780827,https://old.reddit.com/r/Jokes/comments/4pnc9a/breakups_are_hard_britain_should_just_be_like/,self.jokes,,[deleted],Breakups are hard. Britain should just be like,0
post,4pnbes,2qh72,jokes,false,1466780558,https://old.reddit.com/r/Jokes/comments/4pnbes/the_redcoats_are_leaving_the_redcoats_are_leaving/,self.jokes,,[removed],"The Redcoats are leaving, the Redcoats are leaving!",1
post,4pnbc6,2qh72,jokes,false,1466780532,https://old.reddit.com/r/Jokes/comments/4pnbc6/a_jewish_man_sends_his_son_to_israel_to_live/,self.jokes,,"A Jewish man sends his son to Israel to live there for a while. Eventually he returns home and he is now a Christian.  The man finds this to be odd and mentions it to his friend.

The friend listens, thinks for a moment and says, ""That's odd.  I sent my son to Israel as a Jew and he returned as a Christian.""  So the two of them went to see the Rabbi.  

They told the Rabbi the story of how they had both sent their sons to Israel as Jews, and how both sons had returned as Christians.  The Rabbi listened, thought for a minute and then said ""That's odd.  I also sent my son to Israel as a Jew and he returned as a Christian.""

So the three of them decide to go to Israel to find out what's going on over there.  The arrive and go straight to the Western Wall to pray.  They explain to God all about how they sent their sons to Israel as Jews and how the all returned as Christians.""

There is a long silence, and then God begins to speak saying, ""That's odd . . . """,A Jewish man sends his son to Israel to live there for a while . . .,32013
post,4pnbam,2qh72,jokes,false,1466780519,https://old.reddit.com/r/Jokes/comments/4pnbam/whats_the_leading_cause_of_weight_gain_in_women/,self.jokes,,Marriage,What's the leading cause of weight gain in women?,1
post,4pnb8s,2qh72,jokes,false,1466780500,https://old.reddit.com/r/Jokes/comments/4pnb8s/to_be_remain_crowd_in_britain_come_to_canada/,self.jokes,,[deleted],"To be ""Remain"" crowd in Britain... come to Canada!",2
post,4pna5g,2qh72,jokes,false,1466780147,https://old.reddit.com/r/Jokes/comments/4pna5g/why_do_asian_women_have_small_tits/,self.jokes,,Because only A's are acceptable.,Why do Asian women have small tits?,356
post,4pn9ze,2qh72,jokes,false,1466780083,https://old.reddit.com/r/Jokes/comments/4pn9ze/europe_has_freed_up_some_space_today/,self.jokes,,[deleted],Europe has freed up some space today,1
post,4pn9mf,2qh72,jokes,false,1466779962,https://old.reddit.com/r/Jokes/comments/4pn9mf/the_eu_now_has_1_gb_free_space/,self.jokes,,[removed],The EU now has 1 GB free space.,1
post,4pn97e,2qh72,jokes,false,1466779819,https://old.reddit.com/r/Jokes/comments/4pn97e/what_happens_when_frogs_park_illegally/,self.jokes,,[deleted],What happens when frogs park illegally?,3
post,4pn90x,2qh72,jokes,false,1466779757,https://old.reddit.com/r/Jokes/comments/4pn90x/relationships_are_like_fat_girls/,self.jokes,,[deleted],Relationships are like fat girls,3
post,4pn8q2,2qh72,jokes,false,1466779647,https://old.reddit.com/r/Jokes/comments/4pn8q2/i_saw_a_man_staring_at_a_pile_of_poop_on_the/,self.jokes,,"Concerned, I went up to him and asked ""What's the matter?""

""Human. Fecal.""",I saw a man staring at a pile of poop on the street the other day...,1
post,4pn8ok,2qh72,jokes,false,1466779633,https://old.reddit.com/r/Jokes/comments/4pn8ok/todays_newspaper_headlines/,self.jokes,,"The Times: ""PM David Cameron set to resign.""

Daily Mail: ""Tory wanker gets the boot""",Today's newspaper headlines:,0
post,4pn8l8,2qh72,jokes,false,1466779601,https://old.reddit.com/r/Jokes/comments/4pn8l8/weed/,self.jokes,,Nature's way of saying high,Weed.,5
post,4pn8ew,2qh72,jokes,false,1466779543,https://old.reddit.com/r/Jokes/comments/4pn8ew/my_pullout_game_so_strong/,self.jokes,,[deleted],My pullout game so strong ...,1
post,4pn893,2qh72,jokes,false,1466779492,https://old.reddit.com/r/Jokes/comments/4pn893/breakups_are_tough_you_have_to_be_compassionate/,self.jokes,,[deleted],Breakups are tough. You have to be compassionate. Britain should've written a note.,5
post,4pn812,2qh72,jokes,false,1466779415,https://old.reddit.com/r/Jokes/comments/4pn812/what_did_uk_say_to_eu/,self.jokes,,[deleted],What did UK say to EU?,0
post,4pn7bu,2qh72,jokes,false,1466779200,https://old.reddit.com/r/Jokes/comments/4pn7bu/humpty_dumpty_sat_on_a_wall/,self.jokes,,And was shot down by trump border police,Humpty Dumpty sat on a wall.......,1
post,4pn716,2qh72,jokes,false,1466779109,https://old.reddit.com/r/Jokes/comments/4pn716/did_you_hear_that_they_are_banning_orchestral/,self.jokes,,[deleted],Did you hear that they are banning orchestral music from broadcast TV?,3
post,4pn6wt,2qh72,jokes,false,1466779077,https://old.reddit.com/r/Jokes/comments/4pn6wt/kind_of_ironic/,self.jokes,,[removed],Kind of ironic...,1
post,4pn6qw,2qh72,jokes,false,1466779025,https://old.reddit.com/r/Jokes/comments/4pn6qw/with_the_brexit_news_they_say_the_pound_is_failing/,self.jokes,,"They're calling it the ounce, now.","With the brexit news, they say the pound is failing.",9
post,4pn6ke,2qh72,jokes,false,1466778969,https://old.reddit.com/r/Jokes/comments/4pn6ke/breakups_are_tough/,self.jokes,,"You have to be compassionate. Britain should've written a note. 'It's not EU, it's me'.",Breakups are tough.,0
post,4pn66i,2qh72,jokes,false,1466778859,https://old.reddit.com/r/Jokes/comments/4pn66i/when_rorschach_gets_drunk/,self.jokes,,[deleted],When Rorschach gets drunk...,1
post,4pn5vq,2qh72,jokes,false,1466778777,https://old.reddit.com/r/Jokes/comments/4pn5vq/in_the_falsely_attributed_words_of_paul_revere_on/,self.jokes,,[deleted],In the (falsely attributed) words of Paul Revere on this historic occasion,0
post,4pn5mt,2qh72,jokes,false,1466778705,https://old.reddit.com/r/Jokes/comments/4pn5mt/two_drums_and_a_cymbal_roll_down_a_hill/,self.jokes,,ba dum tss,Two drums and a cymbal roll down a hill,1
post,4pn5me,2qh72,jokes,false,1466778702,https://old.reddit.com/r/Jokes/comments/4pn5me/comedy_news_6_24_16/,self.jokes,,"The UK has left the EU. Now if we could only get the BS to leave the GOP and the DEMS!

This congress has really lowered the bar at accomplishing nothing. Before going on break they agreed they won't get a budget done! Paraplegics do more heavy lifting than these jokers!

Forest fires in the West, Floods out East, Heatwave in the Southwest, &amp; the Cubs are in 1st Place. The End is Near!

Over 1 million Americans are now in same sex marriages. In a completely unrelated story Clay Aikens tour is completely sold out!

I went out with a girl who said ""Don't treat me like a date. Treat me like you would your mom"". So I rifled her purse &amp; stole twenty bucks!

Minneapolis has been voted the best place to celebrate July 4th. Worst place; Chicago, the gun fire covers up the rocket blasts! 

A rare near extinct Amazon fish was found in a New Jersey pond. The man who caught it said it was great with tartar sauce! 

I tried Starbucks decaf soda 'Fizzio'. When I saw what it cost I realized it made me 'estupido'! 

On this day in 1997 the Air Force dismissed Roswell's UFO's saying it was just a publicity stunt by mentalist Kreskin.

Today's Inspirational Thought; Until history finally stops repeating itself...man has learned nothing!

Since fundamentalist believe marriage is between a man &amp; a woman, aren't ALL marriages mixed marriages?



",Comedy News 6 24 16,0
post,4pn5hp,2qh72,jokes,false,1466778665,https://old.reddit.com/r/Jokes/comments/4pn5hp/what_does_david_cameron_do_when_he_gets_put_in/,self.jokes,,[deleted],What does David Cameron do when he gets put in charge of something?,0
post,4pn4wd,2qh72,jokes,false,1466778484,https://old.reddit.com/r/Jokes/comments/4pn4wd/britain_is_like_a_man_on_a_toilet/,self.jokes,,It just wanted to get rid of that shit and leave.,Britain is like a man on a toilet...,5
post,4pn4nq,2qh72,jokes,false,1466778396,https://old.reddit.com/r/Jokes/comments/4pn4nq/the_role_of_queen_of_england/,self.jokes,,[deleted],the role of queen of england..,0
post,4pn37m,2qh72,jokes,false,1466777904,https://old.reddit.com/r/Jokes/comments/4pn37m/you_cant_spell_brexit_without/,self.jokes,,[deleted],You can't spell Brexit without...,0
post,4pn2vr,2qh72,jokes,false,1466777795,https://old.reddit.com/r/Jokes/comments/4pn2vr/why_shouldnt_you_have_a_conversation_under_a_tree/,self.jokes,,There may be leavesdropping,Why shouldn't you have a conversation under a tree in the fall?,51
post,4pn2qc,2qh72,jokes,false,1466777745,https://old.reddit.com/r/Jokes/comments/4pn2qc/if_you_punched_a_random_brit_today/,self.jokes,,There would be a 52% chance they deserved it.,If you punched a random Brit today...,3
post,4pn2lp,2qh72,jokes,false,1466777696,https://old.reddit.com/r/Jokes/comments/4pn2lp/what_do_the_mafia_and_a_pussy_have_in_common/,self.jokes,,One slip of the tongue and you're deep in shit.,What do the Mafia and a pussy have in common?,19
post,4pn2l9,2qh72,jokes,false,1466777692,https://old.reddit.com/r/Jokes/comments/4pn2l9/the_brexit_is_obviously_a_result_of_the_uks/,self.jokes,,[deleted],The Brexit is obviously a result of the UK'S strong gun laws...,0
post,4pn2j8,2qh72,jokes,false,1466777673,https://old.reddit.com/r/Jokes/comments/4pn2j8/dj_vu/,self.jokes,,The feeling you get when you've heard the same music in a club before.,DJ vu.,5
post,4pn2hv,2qh72,jokes,false,1466777660,https://old.reddit.com/r/Jokes/comments/4pn2hv/what_happens_when_you_vote_as_a_joke/,self.jokes,,Brexit.,What happens when you vote as a joke?,0
post,4pn2by,2qh72,jokes,false,1466777595,https://old.reddit.com/r/Jokes/comments/4pn2by/eu_just_freed_up_some_space/,self.jokes,,[deleted],EU just freed up some space !,2
post,4pn1zr,2qh72,jokes,false,1466777470,https://old.reddit.com/r/Jokes/comments/4pn1zr/can_i_buy_a_couple_pounds_for_a_dollar/,self.jokes,,[deleted],Can I buy a couple pounds for a dollar?,0
post,4pn0ry,2qh72,jokes,false,1466777039,https://old.reddit.com/r/Jokes/comments/4pn0ry/i_wish_my_girlfriend_went_down_as_much/,self.jokes,,as the pound did last night. ,I wish my girlfriend went down as much...,128
post,4pn0b7,2qh72,jokes,false,1466776875,https://old.reddit.com/r/Jokes/comments/4pn0b7/brexit_to_be_followed_by_grexit_departugal/,self.jokes,,[deleted],Brexit' to be followed by Grexit. De-partugal. Italeave. Fruckoff. Czechout. Oustria. Finish. Slovakout. Latervia. Byegium.,1
post,4pn07g,2qh72,jokes,false,1466776843,https://old.reddit.com/r/Jokes/comments/4pn07g/_/,self.jokes,,[removed],🤔🇪🇺🔚🔜,1
post,4pmzle,2qh72,jokes,false,1466776613,https://old.reddit.com/r/Jokes/comments/4pmzle/what_is_big_black_and_long/,self.jokes,,The lines at KFC,What is big black and long.,38
post,4pmzei,2qh72,jokes,false,1466776541,https://old.reddit.com/r/Jokes/comments/4pmzei/jack_off_all_trades/,self.jokes,,master onan,jack off all trades,0
post,4pmz17,2qh72,jokes,false,1466776410,https://old.reddit.com/r/Jokes/comments/4pmz17/i_feel_quite_light_today/,self.jokes,,Pounds aren't what they used to be.,I feel quite light today.,22
post,4pmyzd,2qh72,jokes,false,1466776391,https://old.reddit.com/r/Jokes/comments/4pmyzd/a_rabbit_and_a_bear/,self.jokes,,"A rabbit and a bear go to relieve themselves in a forest. 
The bear asks the rabbit ""do you have problems with poo sticking you fur?""
""No"" says the rabbit. 
The bear then wipes his bottom with the rabbit. ",A Rabbit and a Bear..,1
post,4pmyqc,2qh72,jokes,false,1466776281,https://old.reddit.com/r/Jokes/comments/4pmyqc/logedy_is_friendly_unless_fed/,self.jokes,,"logedy has been a close friend of mine for a few years, now. yeah, I know, it's a funny name and all, but what can I say? I'm pretty much the same. Quite frankly, logedy sounds like a game of an adventurer who goes by the name of it. specifically, an adventurer of powerful magic -- perhaps even a mage, who's sole destiny is only but to find a magical star that fell onto to earth that is said only to appear everyone one in ten billion years, but contains immense power that if used by a mage, could boost his own power, tenfold!","Logedy is friendly, unless fed.",0
post,4pmynp,2qh72,jokes,false,1466776251,https://old.reddit.com/r/Jokes/comments/4pmynp/britain_do_you/,self.jokes,,[deleted],Britain... do you,0
post,4pmylp,2qh72,jokes,false,1466776234,https://old.reddit.com/r/Jokes/comments/4pmylp/rumour/,self.jokes,,"I heard a rumour that a man in town is selling a fake bedside-clock.

It's a false alarm.",Rumour...,14
post,4pmyf1,2qh72,jokes,false,1466776169,https://old.reddit.com/r/Jokes/comments/4pmyf1/asked_my_coworker_if_saw_the_big_news_report/,self.jokes,,"He said which one, The Mac 'n Cheetos announcement or the UK doing something?


True story, from 3 min ago... 'Murica",Asked my co-worker if saw the big news report...,7
post,4pmyc5,2qh72,jokes,false,1466776139,https://old.reddit.com/r/Jokes/comments/4pmyc5/my_friend_told_me_to_go_to_a_gas_station_cause_he/,self.jokes,,"I told him: ""Urine trouble!""",My friend told me to go to a gas station cause he really had to pee.,0
post,4pmy4v,2qh72,jokes,false,1466776057,https://old.reddit.com/r/Jokes/comments/4pmy4v/gandhi_goes_to_the_barbershop/,self.jokes,,"Gandhi wanted a to get to the barbershop, but he couldn't because there was a river blocking his way. On his side of the river there is a tree and below the tree there are broken branches. On the other side there was a kayak that was just sitting there. Gandhi did not know how to swim so how did he get across the river?
-
-
-
-
-
-
-
-
-
Answer: He didn't because he was bald",Gandhi goes to the barbershop,0
post,4pmy0z,2qh72,jokes,false,1466776011,https://old.reddit.com/r/Jokes/comments/4pmy0z/why_did_the_slave_cross_the_road/,self.jokes,,He didn't have a choice,Why did the slave cross the road?,0
post,4pmxxj,2qh72,jokes,false,1466775969,https://old.reddit.com/r/Jokes/comments/4pmxxj/why_was_6_afraid_of_7/,self.jokes,,[deleted],Why was 6 afraid of 7?,0
post,4pmxgx,2qh72,jokes,false,1466775803,https://old.reddit.com/r/Jokes/comments/4pmxgx/whats_fast_and_can_breathe_underwater/,self.jokes,,"Not a toddler, I can tell you that",What's fast and can breathe underwater?,74
post,4pmx5f,2qh72,jokes,false,1466775687,https://old.reddit.com/r/Jokes/comments/4pmx5f/my_girlfriend_wants_to_go_to_the_uk/,self.jokes,,"I said,""I would rather see EU buy a weightloss program.""",My Girlfriend wants to go to the UK...,0
post,4pmwt9,2qh72,jokes,false,1466775564,https://old.reddit.com/r/Jokes/comments/4pmwt9/nsfw_i_got_an_awesome_handjob_from_my_barber/,self.jokes,,Just one of the many benefits to cutting your own hair,[NSFW] I got an awesome handjob from my barber after my haircut,3
post,4pmw4d,2qh72,jokes,false,1466775313,https://old.reddit.com/r/Jokes/comments/4pmw4d/referendum_results_lead_to_petition_to_stop/,self.jokes,," I mean... uhh... leads to children creating petition because they can't handle the democratic process.*

My mistake!",Referendum results lead to petition to stop children taking part in democratic process...,0
post,4pmw17,2qh72,jokes,false,1466775282,https://old.reddit.com/r/Jokes/comments/4pmw17/i_dont_know_how_valve_managed_to_do_it_but/,self.jokes,,they even included the British Pound in their summer sale this year.,"I don't know how Valve managed to do it, but...",11
post,4pmw01,2qh72,jokes,false,1466775269,https://old.reddit.com/r/Jokes/comments/4pmw01/making_sandwiches_nsfw/,self.jokes,,"A teenage girl wants to take her boyfriend home to have sex, but she shares a bunk bed with her little brother. So they develop code words so the brother won't know what's going on. When she says ""pickles"" he goes faster and when she says ""tomatoes"" he goes slower. 
The next morning the brother asked what she had been doing all night when she tells him ""I was making sandwiches for today's lunch!""
That's when her brother replies, ""oh thank god, i was worried you were fucking your boyfriend but it was just mayonaise on my pillow then last night!""",Making sandwiches (NSFW),1
post,4pmvqy,2qh72,jokes,false,1466775176,https://old.reddit.com/r/Jokes/comments/4pmvqy/please_england_dont_leave/,self.jokes,,[deleted],"Please England, don't leave…",0
post,4pmva4,2qh72,jokes,false,1466775006,https://old.reddit.com/r/Jokes/comments/4pmva4/if_the_leave_camp_was_a_bit_more_subtle_about/,self.jokes,,[deleted],"If the leave camp was a bit more subtle about their victory, it would just be a...",0
post,4pmusl,2qh72,jokes,false,1466774818,https://old.reddit.com/r/Jokes/comments/4pmusl/what_do_you_call_the_dump_you_take_after_a_brunch/,self.jokes,,Brexit.,What do you call the dump you take after a brunch?,0
post,4pmtv3,2qh72,jokes,false,1466774450,https://old.reddit.com/r/Jokes/comments/4pmtv3/what_did_the_electrical_engineer_do_when_she/,self.jokes,,She soldered on. ,What did the electrical engineer do when she found out that she hadn't won the lottery?,1
post,4pmtpj,2qh72,jokes,false,1466774390,https://old.reddit.com/r/Jokes/comments/4pmtpj/where_do_most_black_people_work/,self.jokes,,In jail,Where do most black people work?,0
post,4pmsxb,2qh72,jokes,false,1466774098,https://old.reddit.com/r/Jokes/comments/4pmsxb/what_did_the_eu_get_from_the_uk_leaving_it/,self.jokes,,[deleted],What did the EU get from the UK leaving it?,0
post,4pmsdd,2qh72,jokes,false,1466773861,https://old.reddit.com/r/Jokes/comments/4pmsdd/being_irish_whats_bonos_favorite_song/,self.jokes,,[deleted],"Being irish, Whats Bono's favorite song?",0
post,4pms54,2qh72,jokes,false,1466773775,https://old.reddit.com/r/Jokes/comments/4pms54/my_favorite_rapper_is_50_cent/,self.jokes,,"Or as the British people now call him, 10,000 pounds.",My favorite rapper is 50 cent,1015
post,4pms42,2qh72,jokes,false,1466773761,https://old.reddit.com/r/Jokes/comments/4pms42/the_joke_lies_in_the_comments/,self.jokes,,[removed],The joke lies in the comments.,1
post,4pms1o,2qh72,jokes,false,1466773735,https://old.reddit.com/r/Jokes/comments/4pms1o/after_leaving_the_pm_post_cameron_will_become_a/,self.jokes,,[deleted],"After leaving the PM post, Cameron will become a rapper...",0
post,4pms0r,2qh72,jokes,false,1466773725,https://old.reddit.com/r/Jokes/comments/4pms0r/how_many_brits_are_needed_to_change_a_light_bulb/,self.jokes,,None they just terminate their apartment  contract.,How many brits are needed to change a light bulb,6
post,4pmr83,2qh72,jokes,false,1466773424,https://old.reddit.com/r/Jokes/comments/4pmr83/britain/,self.jokes,,[removed],Britain,1
post,4pmqpl,2qh72,jokes,false,1466773245,https://old.reddit.com/r/Jokes/comments/4pmqpl/a_muslim_terrorist_walks_in_to_a_bar/,self.jokes,,[removed],A Muslim terrorist walks in to a bar..,0
post,4pmqm4,2qh72,jokes,false,1466773208,https://old.reddit.com/r/Jokes/comments/4pmqm4/can_you_remember_the_punch_line_to_that_one/,self.jokes,,Because I lost it.,Can you remember the punch line to that one hilarious joke on here the other day?,0
post,4pmqcc,2qh72,jokes,false,1466773102,https://old.reddit.com/r/Jokes/comments/4pmqcc/what_was_the_cure_for_britains_headache/,self.jokes,,Aleve.,What was the cure for Britain's headache?,0
post,4pmq6t,2qh72,jokes,false,1466773040,https://old.reddit.com/r/Jokes/comments/4pmq6t/brexit_fallout_my_french_toast_has_just/,self.jokes,,and my Irish coffee is drunk.  Again. ,Brexit fallout: my French Toast has just surrendered to my English Muffins. Germany is sending in the Luftwaffle... these events could engulf the entire continental breakfast.,76
post,4pmptj,2qh72,jokes,false,1466772871,https://old.reddit.com/r/Jokes/comments/4pmptj/brexit_related/,self.jokes,,[deleted],Brexit related?,0
post,4pmpo4,2qh72,jokes,false,1466772807,https://old.reddit.com/r/Jokes/comments/4pmpo4/boris_johnson_and_donald_trump_walk_into_a_bar/,self.jokes,,It catches fire. Luckily nothing of value is lost.,Boris Johnson and Donald Trump walk into a bar.,0
post,4pmple,2qh72,jokes,false,1466772777,https://old.reddit.com/r/Jokes/comments/4pmple/european_union/,self.jokes,,THE UK ISN'T IN IT ANYMORE.,EUROPEAN UNION.,0
post,4pmoys,2qh72,jokes,false,1466772527,https://old.reddit.com/r/Jokes/comments/4pmoys/seems_like_a_good_day_to_start_a_diet/,self.jokes,,[deleted],Seems like a good day to start a diet,1
post,4pmovm,2qh72,jokes,false,1466772490,https://old.reddit.com/r/Jokes/comments/4pmovm/song_of_the_day/,self.jokes,,U2: With or without EU,Song of the day:,0
post,4pmoo1,2qh72,jokes,false,1466772413,https://old.reddit.com/r/Jokes/comments/4pmoo1/the_british_pound/,self.jokes,,[removed],The British Pound,1
post,4pmof4,2qh72,jokes,false,1466772302,https://old.reddit.com/r/Jokes/comments/4pmof4/why_was_the_redneck_fired_on_his_first_day/,self.jokes,,[deleted],Why was the redneck fired on his first day manning the missile silo?,0
post,4pmoei,2qh72,jokes,false,1466772291,https://old.reddit.com/r/Jokes/comments/4pmoei/what_did_england_say_to_scotland/,self.jokes,,Send my love to your EU lover,What did England say to Scotland?,0
post,4pmna0,2qh72,jokes,false,1466771795,https://old.reddit.com/r/Jokes/comments/4pmna0/a_happily_married_couple/,self.jokes,,[deleted],A happily married couple....,2
post,4pmn6m,2qh72,jokes,false,1466771761,https://old.reddit.com/r/Jokes/comments/4pmn6m/im_46_and_my_mum_told_me_i_have_to_move_out/,self.jokes,,[deleted],I'm 46 and my Mum told me I have to move out...,0
post,4pmmou,2qh72,jokes,false,1466771551,https://old.reddit.com/r/Jokes/comments/4pmmou/i_regret_joining_the_gym_recently/,self.jokes,,leaving the EU would've been a more effective way to lose pounds ,I regret joining the gym recently..,615
post,4pmmg7,2qh72,jokes,false,1466771452,https://old.reddit.com/r/Jokes/comments/4pmmg7/breaking_europe_awaiting_a_new_wave_of_economical/,self.jokes,,But atleast their English is bloody excellent!,BREAKING: Europe awaiting a new wave of economical refugees!,8
post,4pmm47,2qh72,jokes,false,1466771317,https://old.reddit.com/r/Jokes/comments/4pmm47/nsfw_nsfl_did_you_hear_about_the_the_person_that/,self.jokes,,He rectum.,[NSFW] [NSFL] Did you hear about the the person that made all the butts fall out?,0
post,4pmlle,2qh72,jokes,false,1466771083,https://old.reddit.com/r/Jokes/comments/4pmlle/condoms_prevent_pregnancy/,self.jokes,,and other STDs.,Condoms prevent pregnancy..,1
post,4pml6f,2qh72,jokes,false,1466770889,https://old.reddit.com/r/Jokes/comments/4pml6f/breast_feeding/,self.jokes,,"A blonde woman is walking down the street, with her blouse open. A cop is approaching from about a block away, thinking, ""Boy, my eyes must be going, it looks like that woman's right breast is hanging out."" As he gets closer it becomes apparent that her breast is hanging out. When he gets face to face with her he says, ""Ma'am, are you aware I could cite you for indecent exposure?"" She says, ""Why, officer?"" ""Well, your breast is hanging out."" She looks down and says ""OMIGOD, I left the baby on the bus!"" ",Breast Feeding,12
post,4pmkz9,2qh72,jokes,false,1466770801,https://old.reddit.com/r/Jokes/comments/4pmkz9/so_today_i_woke_up_and_asked_my_uk_counterpart/,self.jokes,,"""Did you have eggs and bacon with your Brexit this morning?""","So, today I woke up and asked my UK counterpart...",0
post,4pmkn1,2qh72,jokes,false,1466770646,https://old.reddit.com/r/Jokes/comments/4pmkn1/does_donald_trump_master_his_tracks/,self.jokes,,Nope. He puts a limiter on there and brick walls it.,Does Donald Trump master his tracks?,1
post,4pmjrk,2qh72,jokes,false,1466770232,https://old.reddit.com/r/Jokes/comments/4pmjrk/eu_referendum/,self.jokes,,"Ok. Bear with me.

All the celebrity deaths in 2016. Missing persons being discussed on Radio 4. Britain votes to leave the EU which leads to David Cameron resigning as PM. The options to replace him include Jeremy Hunt (a deaths eater if ever O saw one). This leads to my conclusion:

Voldemort Has returned! ",EU referendum,0
post,4pmjqs,2qh72,jokes,false,1466770226,https://old.reddit.com/r/Jokes/comments/4pmjqs/todays_friday_so_at_work_im_just_going_to_shoot/,self.jokes,,[removed],"Today's Friday, so at work I'm just going to shoot for amateurductivity.",1
post,4pmjns,2qh72,jokes,false,1466770189,https://old.reddit.com/r/Jokes/comments/4pmjns/the_british_economy/,self.jokes,,[removed],The British Economy,1
post,4pmjga,2qh72,jokes,false,1466770103,https://old.reddit.com/r/Jokes/comments/4pmjga/lets_rename_earth_to_earf_we_need_your_help/,self.jokes,,[removed],Let's Rename Earth to Earf: We Need Your Help!,1
post,4pmjg2,2qh72,jokes,false,1466770102,https://old.reddit.com/r/Jokes/comments/4pmjg2/why_didnt_the_toilet_paper_cross_the_road/,self.jokes,,Because it was stuck in a crack. ,Why didn't the toilet paper cross the road?,5
post,4pmjbr,2qh72,jokes,false,1466770050,https://old.reddit.com/r/Jokes/comments/4pmjbr/what_is_the_capital_of_greece/,self.jokes,,More than the capital of the UK.,What is the capital of Greece?,75
post,4pmj11,2qh72,jokes,false,1466769917,https://old.reddit.com/r/Jokes/comments/4pmj11/whats_a_skydivers_favorite_spice_ground_cumin/,self.jokes,,As long as they aren't running out of thyme.,What's a skydiver's favorite spice? Ground cumin!,2
post,4pmj0b,2qh72,jokes,false,1466769909,https://old.reddit.com/r/Jokes/comments/4pmj0b/a_family_dinner/,self.jokes,,"A family is at the dinner table, when the son asks the father, “Dad, how many kinds of boobs are there?” 

The father, surprised, answers, “Well, son, a woman goes through three phases. In her 20s, a woman’s breasts are like melons, round and firm. In her 30s and 40s, they are like pears, still nice, hanging a bit. After 50, they are like onions.” 

“Onions?” the son asks. 

“Yes. You see them and they make you cry.”

This infuriated his wife and daughter. 

The daughter asks, “Mom, how many different kinds of willies are there?” 

The mother smiles and says, “Well, dear, a man goes through three phases also. In his 20s, his willy is like an oak tree, mighty and hard. In his 30s and 40s, it’s like a birch, flexible but reliable. After his 50s, it’s like a Christmas tree.” 

“A Christmas tree?” the daughter asks.

“Yes, dead from the root up and the balls are just for decoration.”",A family dinner...,47
post,4pmita,2qh72,jokes,false,1466769818,https://old.reddit.com/r/Jokes/comments/4pmita/uk_referendum/,self.jokes,,I hope my grades won't drop as hard as the UK economy. ,UK referendum,0
post,4pmim3,2qh72,jokes,false,1466769736,https://old.reddit.com/r/Jokes/comments/4pmim3/a_man_walks_into_a_bar/,self.jokes,,"A man walks into a bar and sees a beautiful women. He goes over, sits next to her, and gets a drink. After sitting for a minute, he chuckles to himself. 

""What's so funny"" asks the women. 

""I was gonna tell you a joke about my dick but it's too long""

""Oh"" she says "" I'd tell you one about my pussy, but you'll never get it""

",A man walks into a bar...,1
post,4pmihf,2qh72,jokes,false,1466769683,https://old.reddit.com/r/Jokes/comments/4pmihf/i_think_the_uk_shouldve_stayed_in_the_eu/,self.jokes,,But that's just my 2 cents (£12.73),I think the UK should've stayed in the EU.,2
post,4pmie1,2qh72,jokes,false,1466769643,https://old.reddit.com/r/Jokes/comments/4pmie1/what_do_they_say_when_batman_catches_a_cold/,self.jokes,,He's ben affleckted.,What do they say when batman catches a cold?,2
post,4pmibj,2qh72,jokes,false,1466769613,https://old.reddit.com/r/Jokes/comments/4pmibj/a_police_officer_was_interrogating_a_suspect_in_a/,self.jokes,,"""No you see, I couldn't have done it! I was working at the bakery all night making doughnuts!"" ""I'm afraid I'm going to have to place you under arrest. There are too many holes in your story.""",A police officer was interrogating a suspect in a murder case,1
post,4pmia0,2qh72,jokes,false,1466769594,https://old.reddit.com/r/Jokes/comments/4pmia0/i_cant_live_without_eu/,self.jokes,,[deleted],I can't live without EU,0
post,4pmhw7,2qh72,jokes,false,1466769405,https://old.reddit.com/r/Jokes/comments/4pmhw7/what_do_you_call_a_mexican_that_had_his_car_stolen/,self.jokes,,Carloss ,What do you call a Mexican that had his car stolen?,17
post,4pmhr3,2qh72,jokes,false,1466769349,https://old.reddit.com/r/Jokes/comments/4pmhr3/nit_d_kingdom/,self.jokes,,[removed],_nit_d Kingdom,3
post,4pmhot,2qh72,jokes,false,1466769326,https://old.reddit.com/r/Jokes/comments/4pmhot/after_britain_left/,self.jokes,,The EU now has 1GB free,After Britain left...,1
post,4pmhoh,2qh72,jokes,false,1466769322,https://old.reddit.com/r/Jokes/comments/4pmhoh/keep_calm_and/,self.jokes,,PANIC LIKE FUCK!,Keep Calm and,0
post,4pmhlp,2qh72,jokes,false,1466769282,https://old.reddit.com/r/Jokes/comments/4pmhlp/an_egg_voted_to_leave_the_omelet/,self.jokes,,"and then.. it.. did..

yeah, sorry its just too scrambled.

there's no way to get a good yolk out of this mess..",An egg voted to leave the omelet..,1
post,4pmhhk,2qh72,jokes,false,1466769231,https://old.reddit.com/r/Jokes/comments/4pmhhk/theres_some_free_space_in_the_eu_now/,self.jokes,,"1 GB, to be precise.",There's some free space in the EU now..,1
post,4pmg2m,2qh72,jokes,false,1466768586,https://old.reddit.com/r/Jokes/comments/4pmg2m/when_i_lived_in_florida_i_worked_in_an_orange/,self.jokes,,But I got canned for not being able to concentrate,When I lived in Florida I worked in an orange factory..,1
post,4pmfn4,2qh72,jokes,false,1466768382,https://old.reddit.com/r/Jokes/comments/4pmfn4/nsfw_good_luck_mr_collins/,self.jokes,,"Two astronauts successfully landed on the moon and transmitted their thoughts and feelings back to mission control. They described the moon's surface, the atmosphere, the temperature and their feelings of elation at being there. 

Just as the transmission was going off, one of the astronauts was heard to say, ""Good Luck Mr Collins"".

When the men eventually returned to earth, there was lot of media attention but when it came to the meaning of"" Good Luck Mr Collins"", the astronaut refused to explain. 

25 years later, on the anniversary of the moon landing, once again the two astronauts become the centre of attention. It was then, on a late night television programme that the meaning of ""Good Luck Mr Collins"" was explained.

""When I was a young boy, our family lived next door to Mr and Mrs Collins,"" he began, ""and one day, when I was playing in the garden, I heard voices coming from their open bed room window. I heard Mrs Collins yelling at her husband, 

'Oral Sex, that's what you want? Is it... Oral Sex? Let me tell you, when the boy next door lands on moon, then you'll get Oral Sex!' ""","[NSFW] ""Good Luck Mr Collins""",13
post,4pmfk1,2qh72,jokes,false,1466768339,https://old.reddit.com/r/Jokes/comments/4pmfk1/english_man_reaches_for_his_wallet_to_pay_hooker/,self.jokes,,"She replies ""oh, so you want me to pound you?""",English man reaches for his wallet to pay hooker....,1
post,4pmfi6,2qh72,jokes,false,1466768312,https://old.reddit.com/r/Jokes/comments/4pmfi6/why_did_the_pound_crash_after_the_eu_referendum/,self.jokes,,Because the Brexit rexit,Why did the pound crash after the eu referendum?,0
post,4pmfcb,2qh72,jokes,false,1466768231,https://old.reddit.com/r/Jokes/comments/4pmfcb/what_did_uk_say_while_leaving/,self.jokes,,"It's not EU, it's me",What did UK say while leaving?,0
post,4pmf8f,2qh72,jokes,false,1466768175,https://old.reddit.com/r/Jokes/comments/4pmf8f/im_getting_ready_for_lettuce_referendum/,self.jokes,,Leaf or Romaine.,I'm getting ready for Lettuce Referendum...,0
post,4pmevk,2qh72,jokes,false,1466768007,https://old.reddit.com/r/Jokes/comments/4pmevk/an_englishman_an_irishman_a_welshman_and_a/,self.jokes,,Then a few decades later they walk out again squabbling among themselves.,"An Englishman, an Irishman, a Welshman, and a Scotsman walk into a bar.",2
post,4pmdx6,2qh72,jokes,false,1466767501,https://old.reddit.com/r/Jokes/comments/4pmdx6/a_salesman_knocks_on_the_door_of_a_house/,self.jokes,,"It is opened by a young girl, maybe 12 or 13. She is heavily made up, her hair is dyed and permed, and she is dressed in a short skirt and a low-cut top. In one hand, she holds a cigarette holder, in the other a glass of whisky. Behind her, the salesman sees two naked men in bondage gear.

""Er...hello Miss"", he says cautiously. ""Are your parents home?""

The girl just looks at him. ""What do you think?""",A salesman knocks on the door of a house...,1
post,4pmdgs,2qh72,jokes,false,1466767262,https://old.reddit.com/r/Jokes/comments/4pmdgs/want_to_hear_a_racist_joke/,self.jokes,,[removed],Want to hear a racist joke?,4
post,4pmdev,2qh72,jokes,false,1466767236,https://old.reddit.com/r/Jokes/comments/4pmdev/the_uk_could_be_the_51st_state/,self.jokes,,It'd just be like moving in with your grandson. ,The UK could be the 51st State.,4
post,4pmddc,2qh72,jokes,false,1466767212,https://old.reddit.com/r/Jokes/comments/4pmddc/bacon_may_cause_cancer/,self.jokes,,[deleted],"""Bacon may cause cancer...""",0
post,4pmdcb,2qh72,jokes,false,1466767198,https://old.reddit.com/r/Jokes/comments/4pmdcb/a_muslim_walks_into_a_bar_and_the_bartender_asks/,self.jokes,,[removed],"A Muslim walks into a bar and the bartender asks ""what'll you have""?",0
post,4pmd17,2qh72,jokes,false,1466767049,https://old.reddit.com/r/Jokes/comments/4pmd17/how_much_space_did_the_eu_gain/,self.jokes,,[removed],How much space did the EU gain?,0
post,4pmcwa,2qh72,jokes,false,1466766972,https://old.reddit.com/r/Jokes/comments/4pmcwa/i_was_walking_in_the_countryside/,self.jokes,,I asked a wind generator what kind of music it liked. It was a big metal fan.,I was walking in the countryside.,1
post,4pmcew,2qh72,jokes,false,1466766740,https://old.reddit.com/r/Jokes/comments/4pmcew/i_can_only_get_off_to_numbers_now/,self.jokes,,[deleted],I can only get off to numbers now.,2
post,4pmbhn,2qh72,jokes,false,1466766279,https://old.reddit.com/r/Jokes/comments/4pmbhn/nigel_farage_isnt_too_happy_about_the_result_of/,self.jokes,,Leave won by a minority.,Nigel Farage isn't too happy about the result of the EU Referendum.,1
post,4pmbgl,2qh72,jokes,false,1466766263,https://old.reddit.com/r/Jokes/comments/4pmbgl/and_then_the_brit_said/,self.jokes,,[deleted],And then the Brit said...,6
post,4pmasy,2qh72,jokes,false,1466765915,https://old.reddit.com/r/Jokes/comments/4pmasy/how_will_the_eu_die/,self.jokes,,[deleted],How will the EU die?,1
post,4pmarj,2qh72,jokes,false,1466765892,https://old.reddit.com/r/Jokes/comments/4pmarj/so_the_uk_voted_to_leave_the_eu_today/,self.jokes,,[removed],So the UK voted to leave the EU today...,1
post,4pmam6,2qh72,jokes,false,1466765817,https://old.reddit.com/r/Jokes/comments/4pmam6/so_a_duck_walks_into_a_pharmacy/,self.jokes,,and says “Give me some chap-stick… and put it on my bill.,So a duck walks into a pharmacy,1
post,4pmajo,2qh72,jokes,false,1466765777,https://old.reddit.com/r/Jokes/comments/4pmajo/the_uk_will_go_blind/,self.jokes,,Too much playing with your Johnson does that.,The UK will go blind.,0
post,4pma8h,2qh72,jokes,false,1466765624,https://old.reddit.com/r/Jokes/comments/4pma8h/what_did_the_obstinate_yogi_say_when_asked_to/,self.jokes,,Nah imma stay,What did the obstinate yogi say when asked to leave?,1
post,4pma6i,2qh72,jokes,false,1466765594,https://old.reddit.com/r/Jokes/comments/4pma6i/whats_fun_for_910_people/,self.jokes,,gang-rape,Whats fun for 9/10 people?,7
post,4pm9wu,2qh72,jokes,false,1466765470,https://old.reddit.com/r/Jokes/comments/4pm9wu/my_girlfriend_left_me/,self.jokes,,[removed],My girlfriend left me,1
post,4pm9qu,2qh72,jokes,false,1466765385,https://old.reddit.com/r/Jokes/comments/4pm9qu/what_did_the_frog_say_to_the_hooker/,self.jokes,,"""Stribbit"".

Don't worry fellas, I know my way out.",What did the frog say to the hooker?,0
post,4pm9q8,2qh72,jokes,false,1466765377,https://old.reddit.com/r/Jokes/comments/4pm9q8/britain_no_more_fish_n_chips_for_you/,self.jokes,,[removed],"Britain, no more Fish n' Chips for you",1
post,4pm9l1,2qh72,jokes,false,1466765298,https://old.reddit.com/r/Jokes/comments/4pm9l1/when_someone_asks_if_im_going_out_after_work/,self.jokes,,"Yea, out the door to go home.",When someone asks if I'm going out after work,0
post,4pm9gf,2qh72,jokes,false,1466765234,https://old.reddit.com/r/Jokes/comments/4pm9gf/i_decided_to_go_horseback_riding_yesterday/,self.jokes,,Yesterday was not a good day. I decided to go horseback riding something I haven't done in over 20 years. It turned out to be a big mistake! I got on the horse and started out slow but then we went a little faster and before I knew it we were going as fast as the horse could go. I couldn't take the pace and fell off but caught my foot in the stirrup with the horse dragging me. It wouldn't stop it just kept going around and around in a circle.Thank goodness the store manager at Wal-Mart came out and unplugged the machine.,I decided to go horseback riding yesterday,1
post,4pm9er,2qh72,jokes,false,1466765207,https://old.reddit.com/r/Jokes/comments/4pm9er/you_really_have_to_admire_brits_who_voted_to_leave/,self.jokes,,They were so worried about immigrants ruining their economy than they preempted it by doing it themselves.,you really have to admire brits who voted to leave,90
post,4pm8qq,2qh72,jokes,false,1466764865,https://old.reddit.com/r/Jokes/comments/4pm8qq/its_important_to_just_accept_the_result_and_move/,self.jokes,,"#...possibly to another country.""

_Frankie Boyle, (Scottish Comedian)_","""It's important to just accept the result and move on",1
post,4pm8o7,2qh72,jokes,false,1466764830,https://old.reddit.com/r/Jokes/comments/4pm8o7/my_mother_caught_me_wanking/,self.jokes,,[deleted],My mother caught me wanking...,0
post,4pm8if,2qh72,jokes,false,1466764750,https://old.reddit.com/r/Jokes/comments/4pm8if/whats_the_worst_thing_to_forget_when_you_post_a/,self.jokes,,[removed],What's the worst thing to forget when you post a joke?,1
post,4pm8gp,2qh72,jokes,false,1466764722,https://old.reddit.com/r/Jokes/comments/4pm8gp/what_do_boris_johnson_the_british_economy_and_an/,self.jokes,,They're all laughing stocks.,"What do Boris Johnson, the British Economy, and an entertained cube of beef extract have in common?",1
post,4pm8fx,2qh72,jokes,false,1466764709,https://old.reddit.com/r/Jokes/comments/4pm8fx/a_snake_walks_into_a_crowded_bar/,self.jokes,,[removed],A snake walks into a crowded bar,1
post,4pm7dc,2qh72,jokes,false,1466764165,https://old.reddit.com/r/Jokes/comments/4pm7dc/you_make_tea_of_every_spices/,self.jokes,,Here is some salttea. ,You make tea of every spices..,0
post,4pm70l,2qh72,jokes,false,1466763983,https://old.reddit.com/r/Jokes/comments/4pm70l/what_is_aquamans_special_ability/,self.jokes,,[deleted],What is Aquaman's special ability?,0
post,4pm6gv,2qh72,jokes,false,1466763702,https://old.reddit.com/r/Jokes/comments/4pm6gv/how_do_you_become_a_millionaire_in_postbrexit_uk/,self.jokes,,"First, start off with a billion pounds.. ",How do you become a millionaire in post-Brexit UK?,0
post,4pm5o8,2qh72,jokes,false,1466763277,https://old.reddit.com/r/Jokes/comments/4pm5o8/britain_has_a_new_national_anthem/,self.jokes,,[removed],Britain has a new national anthem,1
post,4pm5fs,2qh72,jokes,false,1466763159,https://old.reddit.com/r/Jokes/comments/4pm5fs/gotta_hand_it_to_gay_porn_starts/,self.jokes,,[deleted],Gotta hand it to gay porn starts...,1
post,4pm4w5,2qh72,jokes,false,1466762873,https://old.reddit.com/r/Jokes/comments/4pm4w5/want_to_hear_a_fat_joke/,self.jokes,,[deleted],Want to hear a fat joke?,0
post,4pm4m6,2qh72,jokes,false,1466762729,https://old.reddit.com/r/Jokes/comments/4pm4m6/meanwhile_in_glasgie/,self.jokes,,"People are panic buying nail polish, shoe polish, and even furniture polish.

There seems to have been a wee misunderstanding about which polish won't be in the UK soon.",Meanwhile in Glasgie,1
post,4pm4f5,2qh72,jokes,false,1466762627,https://old.reddit.com/r/Jokes/comments/4pm4f5/how_do_you_call_niggeria_leaving_eu/,self.jokes,,blackout,How do you call Niggeria leaving EU?,0
post,4pm490,2qh72,jokes,false,1466762545,https://old.reddit.com/r/Jokes/comments/4pm490/they_said_brexit_would_let_us_get_closer_to_noneu/,self.jokes,,"They were right, we now have more in common with Zimbabwe than ever before.",They said Brexit would let us get closer to non-EU countries.,29
post,4pm48i,2qh72,jokes,false,1466762534,https://old.reddit.com/r/Jokes/comments/4pm48i/with_the_way_brexit_is_looking_the_pound_will/,self.jokes,,[removed],"With the way Brexit is looking, the Pound will soon become the gram.",1
post,4pm3if,2qh72,jokes,false,1466762129,https://old.reddit.com/r/Jokes/comments/4pm3if/what_do_you_call_it_when_someone_asks_their/,self.jokes,,Scotland.,What do you call it when someone asks their friend to stayas a wingman at a party with them and then sneaks out the backdoor themselves five minutes later?,3
post,4pm376,2qh72,jokes,false,1466761936,https://old.reddit.com/r/Jokes/comments/4pm376/led_zeppelin_predicted_the_brexit/,self.jokes,,"Baby I'm gonna Leave EU

Leave EU when the summer comes

Leave EU when the summer comes a-rolling.",Led Zeppelin predicted the Brexit!,4
post,4pm2ei,2qh72,jokes,false,1466761516,https://old.reddit.com/r/Jokes/comments/4pm2ei/edgy_joke_what_do_you_call_a_guy_who_does/,self.jokes,,The Edge.,Edgy joke: What do you call a guy who does everything pro bono?,1
post,4pm2aw,2qh72,jokes,false,1466761465,https://old.reddit.com/r/Jokes/comments/4pm2aw/hey_wanna_hear_a_joke/,self.jokes,,[deleted],Hey wanna hear a joke,0
post,4pm1mb,2qh72,jokes,false,1466761090,https://old.reddit.com/r/Jokes/comments/4pm1mb/if_jesus_died_for_our_sin/,self.jokes,,Who died for our cos and tan?,if jesus died for our sin...,281
post,4pm0jl,2qh72,jokes,false,1466760480,https://old.reddit.com/r/Jokes/comments/4pm0jl/what_do_we_say_to_boris_johnson_and_donald_trump/,self.jokes,,Hair Hair!,What do we say to Boris Johnson and Donald Trump running the world?,9
post,4pm093,2qh72,jokes,false,1466760316,https://old.reddit.com/r/Jokes/comments/4pm093/my_penis_is_only_three_inches/,self.jokes,,Since that fucker kicked my sisters chin. ,My penis is only three inches...,0
post,4plzvk,2qh72,jokes,false,1466760091,https://old.reddit.com/r/Jokes/comments/4plzvk/cameron/,self.jokes,,Cameroff,Cameron,15
post,4plzql,2qh72,jokes,false,1466760006,https://old.reddit.com/r/Jokes/comments/4plzql/brexit_vote_goes_down_as_one_of_the_brits_most/,self.jokes,,Jarvis Cocker stage invasion during Michael Jackson's 'Earth Song' falls to #2.,Brexit Vote goes down as one of the Brit's most shocking moments...,1
post,4plzki,2qh72,jokes,false,1466759922,https://old.reddit.com/r/Jokes/comments/4plzki/walking_didgeridoo/,self.jokes,,I heard what sounded like a didgeridoo coming down the street one very very windy day. Turns out it was just Michelle Duggar wearing a skirt.,Walking didgeridoo,1
post,4plzfz,2qh72,jokes,false,1466759853,https://old.reddit.com/r/Jokes/comments/4plzfz/how_does_the_uk_commit_suicide/,self.jokes,,[deleted],How does the UK commit suicide?,2
post,4plzb3,2qh72,jokes,false,1466759772,https://old.reddit.com/r/Jokes/comments/4plzb3/i_was_dropped_on_my_head_as_a_baby/,self.jokes,,but not as hard as the pound just dropped. ,I was dropped on my head as a baby,4
post,4plz7l,2qh72,jokes,false,1466759712,https://old.reddit.com/r/Jokes/comments/4plz7l/a_zoophile_a_necrophiliac_a_hunter_and_a_masochist/,self.jokes,,"A zoophile, a necrophiliac, a hunter and a masochist get together in a group.

The hunter says: Alright, the zoophile, you fuck a dog, okay?

The zoophile agrees. The hunter says: ""Then I shoot it, okay? Then the necrophiliac fucks the dog, which is now dead, is that cool?

The necrophiliac agrees. The hunter then says: ""And you, masochist, what would you like to do?"" to which the masochist replies: ""Woof.""","A zoophile, a necrophiliac, a hunter and a masochist...",5
post,4plz5y,2qh72,jokes,false,1466759693,https://old.reddit.com/r/Jokes/comments/4plz5y/now_that_brexit_has_won/,self.jokes,,[deleted],Now that Brexit has won...,0
post,4plz32,2qh72,jokes,false,1466759647,https://old.reddit.com/r/Jokes/comments/4plz32/did_opinion_hear_about_the_european_data_theft/,self.jokes,,They are 1GB short ,Did opinion hear about the European data theft?,0
post,4plz0k,2qh72,jokes,false,1466759602,https://old.reddit.com/r/Jokes/comments/4plz0k/i_saw_an_ad_about_this_tractor_which_wheels_can/,self.jokes,,I guess you can call it a..  pro  tractor,I saw an ad about this tractor which wheels can spin 180 degrees without it moving.,1
post,4plyu0,2qh72,jokes,false,1466759485,https://old.reddit.com/r/Jokes/comments/4plyu0/know_what_i_call_girls_who_run_faster_than_me/,self.jokes,,Cardio  ,Know what I call girls who run faster than me?,2
post,4plyk4,2qh72,jokes,false,1466759310,https://old.reddit.com/r/Jokes/comments/4plyk4/with_britain_voting_to_leave_the_eu_has_lost_some/,self.jokes,,[deleted],"With Britain voting to leave, the EU has lost some space...",1
post,4plyfp,2qh72,jokes,false,1466759240,https://old.reddit.com/r/Jokes/comments/4plyfp/the_us_is_waking_up_to_news_of_brexit_vote_leave/,self.jokes,,Bill Clinton leads 'BJ for Prime Minister' calls.,The US is waking up to news of Brexit 'Vote Leave' win...,4
post,4plxx8,2qh72,jokes,false,1466758946,https://old.reddit.com/r/Jokes/comments/4plxx8/whos_the_rapper_with_the_ability_to_dis_everyone/,self.jokes,,[deleted],Who's the rapper with the ability to dis everyone?,2
post,4plxe7,2qh72,jokes,false,1466758649,https://old.reddit.com/r/Jokes/comments/4plxe7/several_eu_countries_have_also_decided_to_have/,self.jokes,,Grexit. Departugal. Italeave. Fruckoff. Czechout. Oustria. Finish. Slovakout. Latervia. Byegium,Several EU countries have also decided to have referenda on their EU membership. This is what they're called!,1
post,4plx80,2qh72,jokes,false,1466758553,https://old.reddit.com/r/Jokes/comments/4plx80/english_within_the_eu_after_todays_vote/,self.jokes,,"Due to todays vote, The European Commission has announced an agreement whereby English will still remain the official language of the EU, rather than German. Her Majesty's Government conceded that English spelling had room for improvement and has therefore accepted a five-year phasing in of ""Euro-English"".
In the first year, ""s"" will replace the soft ""c"". Sertainly, this will make sivil servants jump for joy. The hard ""c"" will be dropped in favour of the ""k"", Which should klear up some konfusion and allow one key less on keyboards.
There will be growing publik enthusiasm in the sekond year, when the troublesome ""ph"" will be replaced with ""f"", making words like ""fotograf"" 20% shorter.
In the third year, publik akseptanse of the new spelling kan be expekted to reach the stage where more komplikated changes are possible. Governments will enkourage the removal of double letters which have always ben a deterent to akurate speling. Also, al wil agre that the horible mes of the silent ""e"" is disgrasful.
By the fourth yer, peopl wil be reseptiv to steps such as replasing ""th"" with ""z"" and ""w"" with ""v"".
During ze fifz yer, ze unesesary ""o"" kan be dropd from vords kontaining ""ou"" and similar changes vud of kors be aplid to ozer kombinations of leters. After zis fifz yer, ve vil hav a reli sensibl riten styl. Zer vil be no mor trubls or difikultis and everivun vil find it ezi to understand ech ozer. ZE DREM VIL FINALI COM TRU!
Herr Schmidt",English within the EU after todays Vote,0
post,4plwy1,2qh72,jokes,false,1466758366,https://old.reddit.com/r/Jokes/comments/4plwy1/america_is_like_an_insideout_oreo/,self.jokes,,[deleted],America is like an inside-out Oreo.,7
post,4plwdt,2qh72,jokes,false,1466758055,https://old.reddit.com/r/Jokes/comments/4plwdt/the_one_thing_i_hate_about_cliffhangers_is/,self.jokes,,[removed],The one thing I hate about cliffhangers is...,1
post,4plwd1,2qh72,jokes,false,1466758045,https://old.reddit.com/r/Jokes/comments/4plwd1/me_and_the_wife_88ed_last_night/,self.jokes,,"It's like 69'ing, but for fat people.",Me and the wife 88'ed last night.,61
post,4plvu3,2qh72,jokes,false,1466757733,https://old.reddit.com/r/Jokes/comments/4plvu3/never_trust_a_parasol/,self.jokes,,I hear they can be shady.,Never trust a Parasol...,2
post,4plvjf,2qh72,jokes,false,1466757565,https://old.reddit.com/r/Jokes/comments/4plvjf/does_this_mean_that_iceland_automatically_qualify/,self.jokes,,[removed],Does this mean that Iceland automatically qualify?,1
post,4plvbx,2qh72,jokes,false,1466757432,https://old.reddit.com/r/Jokes/comments/4plvbx/the_david_cameron_diet/,self.jokes,,You'll never lose your pounds quicker.,The David Cameron diet:,436
post,4plusi,2qh72,jokes,false,1466757106,https://old.reddit.com/r/Jokes/comments/4plusi/whats_the_difference_between_your_pc_and_your/,self.jokes,,"Usually its small, used often and you dont let just ANYONE touch it.",What's the difference between your PC and your Penis?,0
post,4pluqv,2qh72,jokes,false,1466757086,https://old.reddit.com/r/Jokes/comments/4pluqv/santa_is_never_lonely/,self.jokes,,He has many deer friends,Santa is never lonely,11
post,4plup8,2qh72,jokes,false,1466757063,https://old.reddit.com/r/Jokes/comments/4plup8/britain_just_left_the_eu_but_theyll_be_alright/,self.jokes,,"After all, you always lose a few pounds after a break up.",Britain just left the EU! But they'll be alright...,0
post,4pluoo,2qh72,jokes,false,1466757055,https://old.reddit.com/r/Jokes/comments/4pluoo/i_fucked_myself_last_night/,self.jokes,,I wanted to get first-hand experience.,I fucked myself last night.,24
post,4plu8y,2qh72,jokes,false,1466756775,https://old.reddit.com/r/Jokes/comments/4plu8y/the_one_thing_i_hate_about_cliffhangers_is/,self.jokes,,[removed],The one thing I hate about cliffhangers is...,1
post,4plu0a,2qh72,jokes,false,1466756621,https://old.reddit.com/r/Jokes/comments/4plu0a/europe_be_like/,self.jokes,,"eu: uk bro?

uk: it's not eu, it's me.",Europe be like...,312
post,4pltsv,2qh72,jokes,false,1466756497,https://old.reddit.com/r/Jokes/comments/4pltsv/why_your_girlfriend_is_with_you/,self.jokes,,Because she can't have Rick Malabri. ,Why your girlfriend is with you.,0
post,4pltqw,2qh72,jokes,false,1466756466,https://old.reddit.com/r/Jokes/comments/4pltqw/found_a_shop_store_called_dicks_vape/,self.jokes,,[removed],found a shop store called Dick's Vape,1
post,4pltp8,2qh72,jokes,false,1466756447,https://old.reddit.com/r/Jokes/comments/4pltp8/the_good_news_is_that_i_placed_a_safety_bet_on/,self.jokes,,the bad news is my winnings are in pound sterling.,The good news is that I placed a safety bet on Brexit...,2
post,4pltp0,2qh72,jokes,false,1466756443,https://old.reddit.com/r/Jokes/comments/4pltp0/it_seems_that_theres_a_lot_of_eu_jokes_lately_let/,self.jokes,,[deleted],"It seems that there's a lot of EU jokes lately, let me tell a different one",0
post,4pltgo,2qh72,jokes,false,1466756319,https://old.reddit.com/r/Jokes/comments/4pltgo/a_trip_to_israel/,self.jokes,,[deleted],A Trip to Israel..,1
post,4plt79,2qh72,jokes,false,1466756176,https://old.reddit.com/r/Jokes/comments/4plt79/boy_or_girl/,self.jokes,,"A: Just look at that young person with the short hair and blue jeans. Is it a boy or a girl?
B: It's a girl. She's my daughter.
A: Oh, I'm sorry, sir. I didn't know that you were her father.
B: I'm not. I'm her mother.",Boy or Girl,4
post,4plt5e,2qh72,jokes,false,1466756146,https://old.reddit.com/r/Jokes/comments/4plt5e/the_british_pound/,self.jokes,,You mean the British Ounce.,The British Pound?,3
post,4plsxs,2qh72,jokes,false,1466756021,https://old.reddit.com/r/Jokes/comments/4plsxs/_/,self.jokes,,Vegans,.,0
post,4plsxc,2qh72,jokes,false,1466756016,https://old.reddit.com/r/Jokes/comments/4plsxc/late_one_night_han_and_leia_are_hanging_out/,self.jokes,,"when Leia starts bitching about never being able to understand Chewy. Han, fed up with Leia's attitude replied.....

""look princess, there's nothing I can do about it, that's just the way the wookie mumbles""","Late one night, Han and Leia are hanging out getting a bit drunk....",102
post,4plsrn,2qh72,jokes,false,1466755915,https://old.reddit.com/r/Jokes/comments/4plsrn/what_do_eskimos_and_tupperware_have_in_common/,self.jokes,,They both love a tight seal! ,What do Eskimos and Tupperware have in common?,11
post,4plskx,2qh72,jokes,false,1466755805,https://old.reddit.com/r/Jokes/comments/4plskx/i_wanted_to_tell_a_gay_joke_in_light_of_the/,self.jokes,,[deleted],I wanted to tell a gay joke in light of the recent mass shooting...,0
post,4plrw8,2qh72,jokes,false,1466755418,https://old.reddit.com/r/Jokes/comments/4plrw8/good_thing_is_that_the_irish_wont_be_leaving_eu/,self.jokes,," Although, U2 would probably still sound as good With or Without EU.",Good thing is that the Irish won't be leaving EU.,1
post,4plrus,2qh72,jokes,false,1466755395,https://old.reddit.com/r/Jokes/comments/4plrus/living_in_britain/,self.jokes,,[removed],Living in britain,1
post,4plrru,2qh72,jokes,false,1466755350,https://old.reddit.com/r/Jokes/comments/4plrru/whats_the_most_awkward_moment_for_jesus_during_sex/,self.jokes,,When they scream his fathers name.,What's the most awkward moment for Jesus during sex?,3
post,4plrpr,2qh72,jokes,false,1466755311,https://old.reddit.com/r/Jokes/comments/4plrpr/what_do_you_call_a_canadian_and_a_paedophile/,self.jokes,,Alien vs Predator,What do you call a Canadian and a paedophile fighting?,0
post,4pl