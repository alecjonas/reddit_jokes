self.jokes,,Mr. Tyson,What was Mike Tyson's nickname in Prison?,2
post,3kb3mx,2qh72,jokes,false,1441837493,https://old.reddit.com/r/Jokes/comments/3kb3mx/a_brunette_red_head_and_blonde_are_pregnant/,self.jokes,,"A blonde, brunette, and redhead go to the doctor and find out that they are pregnant so they want to find out the sex of the baby. The brunette says, well I was on the bottom so I'm having a boy. The redhead said I was on top so I'm having a girl. The Blonde said, I guess im having puppies!
","A brunette, red head and blonde are pregnant.",8
post,3kb3jw,2qh72,jokes,false,1441837465,https://old.reddit.com/r/Jokes/comments/3kb3jw/an_elderly_couple_decide_to_go_to_the_doctor/,self.jokes,,[deleted],An elderly couple decide to go to the doctor...,8
post,3kb3iz,2qh72,jokes,false,1441837457,https://old.reddit.com/r/Jokes/comments/3kb3iz/blonde_alumna/,self.jokes,,[deleted],Blonde alumna,0
post,3kb3ax,2qh72,jokes,false,1441837373,https://old.reddit.com/r/Jokes/comments/3kb3ax/a_man_is_at_a_party_with_a_bunch_of_his_coworkers/,self.jokes,,"After a couple of hours he's completely wasted. At some point, not knowing what he's doing, the man begins to urinate all over his boss. The man wakes up the next morning with a splitting head ache and no idea what happened the night before. His wife comes up to him and says, ""Bad news, you peed on your boss last night and he fired you."" ""Damn! Well screw him!,"" the man replies. The wife pauses for a second and then says, ""I did, you're back to work on Monday.""",A man is at a party with a bunch of his coworkers and his boss.,4
post,3kb37w,2qh72,jokes,false,1441837342,https://old.reddit.com/r/Jokes/comments/3kb37w/another_little_johnny_joke/,self.jokes,,"On the last day of kindergarten, all the children brought presents for their teacher.  The florist's son handed the teacher a gift.  She shook it, held it up and said, ""I bet I know what it is - it's some flowers!""  ""That's right!"" shouted the little boy.  Then the candy store owner's daughter handed the teacher a gift.  She held it up, shook it and said. ""I bet I know what it is - it's a box of candy!""  ""That's right!"" shouted the little girl.  The next gift was from the liquor store owner's son, Little Johnny.  The teacher held it up and saw that it was leaking.  She touched a drop with her finger and tasted it.  ""Is it wine?"" she asked. ""No,"" Little Johnny answered.  The teacher touched another drop to her tongue. ""Is it champagne?"" she asked.  ""No,"" he answered.  Finally, the teacher said, ""I give up. What is it?""  Little Johnny replied, ""A puppy!""",Another Little Johnny joke,2
post,3kb34x,2qh72,jokes,false,1441837306,https://old.reddit.com/r/Jokes/comments/3kb34x/50_cent_dr_dre_and_eminem_walk_into_a_grocery/,self.jokes,,"Eminem grabs a soda, pays for it at the counter and leaves. 50 cent asks for a pack of swishers, pays for it and leaves. 
""Wait!!!"" screams the clerk as they leave.
Not knowing the man, the two rappers share a confused look and ask him what the problem is.
The clerk sighs and says, ""Come on guys. You Forgot About Dre.""


*****so lame I know, but I haven't seen a rapper joke in a while so.... ","50 Cent, Dr. Dre, and Eminem walk into a grocery store late at night.",1
post,3kb25o,2qh72,jokes,false,1441836968,https://old.reddit.com/r/Jokes/comments/3kb25o/told_my_friends_i_was_taking_my_wife_to_the/,self.jokes,,"One of them said ""Jamaica?""

I said ""No, she wanted to go""",Told my friends I was taking my wife to the Caribbean for our honeymoon,1
post,3kb1dn,2qh72,jokes,false,1441836717,https://old.reddit.com/r/Jokes/comments/3kb1dn/whats_and_electricians_favourite_band/,self.jokes,,AC/DC,What's and electricians favourite band?,0
post,3kb16s,2qh72,jokes,false,1441836651,https://old.reddit.com/r/Jokes/comments/3kb16s/what_do_you_call_a_lesbian_dinosaur/,self.jokes,,Licktalottapuss.,What do you call a lesbian dinosaur.,7
post,3kb14s,2qh72,jokes,false,1441836636,https://old.reddit.com/r/Jokes/comments/3kb14s/what_do_you_call_an_asian_gold_digger/,self.jokes,,Cha Ching,What do you call an Asian gold digger?,79
post,3kb0h4,2qh72,jokes,false,1441836396,https://old.reddit.com/r/Jokes/comments/3kb0h4/how_many_apple_enthusiasts_does_it_take_to_screw/,self.jokes,,[deleted],How many Apple enthusiasts does it take to screw in an Apple brand lightbulb?,0
post,3kb09o,2qh72,jokes,false,1441836326,https://old.reddit.com/r/Jokes/comments/3kb09o/how_do_you_stop_an_italian_from_talking/,self.jokes,,[deleted],How do you stop an Italian from talking?,1
post,3kazpt,2qh72,jokes,false,1441836134,https://old.reddit.com/r/Jokes/comments/3kazpt/i_see_you_7yearold_joke_and_raise_you_mine_why/,self.jokes,,[deleted],I see you 7-year-old joke... And raise you mine: Why are Transformers' (the robots) mother and father never seen in the cartoons?,1
post,3kazoq,2qh72,jokes,false,1441836124,https://old.reddit.com/r/Jokes/comments/3kazoq/little_johnnys_at_it_again/,self.jokes,,"A teacher asks her class, ""What do you want to be when you grow up?"" Little Johnny says ""I wanna be a billionaire, going to the most expensive clubs, take the best bitch with me, give her a Ferrari worth over a million bucks, an apartment in Hawaii, a mansion in Paris, a jet to travel through Europe, an Infinite Visa Card and to make love to her three times a day"". The teacher, shocked, and not knowing what to do with the bad behavior of the child, decides not to give importance to what he said and then continues the lesson. ""And you, Susie? "" the teacher asks. Susie says ""I wanna be Johnny's bitch.""",Little Johnny's at it again....,7
post,3kaz2m,2qh72,jokes,false,1441835898,https://old.reddit.com/r/Jokes/comments/3kaz2m/california/,self.jokes,,"Q: How many Northern Californians does it take to screw in a lightbulb?

A: Hella.",California,15
post,3kayui,2qh72,jokes,false,1441835821,https://old.reddit.com/r/Jokes/comments/3kayui/a_woman_was_in_bed_with_her_lover_when_she_heard/,self.jokes,,"""Hurry!"" she said.  ""Stand in the corner.""  She quickly rubbed baby oil all over him and then she dusted him with talcum powder.  ""Don't move until I tell you to,"" she whispered.  ""Just pretend you're a statue.""

""What's this, honey?"" the husband inquired as he entered the room.

""Oh, it's just a statue,"" she replied nonchalantly.  ""The Smiths bought one for their bedroom.  I liked it so much, I got one for us, too.""

No more was said about the statue, not even later that night when they went to sleep.  

Around two in the morning the husband got out of bed, went to the kitchen and returned a while later with a sandwich and a glass of milk. 

""Here,"" he said to the 'statue'.  ""Eat something.  I stood like an idiot at the Smiths' for three days and nobody offered me as much as a glass of water.""",A woman was in bed with her lover when she heard her husband opening the front door.,7587
post,3kaxj7,2qh72,jokes,false,1441835370,https://old.reddit.com/r/Jokes/comments/3kaxj7/who_is_a_home_repairmans_favorite_rapper/,self.jokes,,[deleted],Who is a home repairman's favorite rapper?,1
post,3kaxed,2qh72,jokes,false,1441835325,https://old.reddit.com/r/Jokes/comments/3kaxed/there_are_only_two_kinds_of_people_in_this_world/,self.jokes,,"Those who pee in the shower, and liars. ",There are only two kinds of people in this world.,1
post,3kaxcs,2qh72,jokes,false,1441835306,https://old.reddit.com/r/Jokes/comments/3kaxcs/have_you_heard_of_the_two_mexican_firemen/,self.jokes,,Hose-A and Hose-B.,Have you heard of the two Mexican firemen?,3
post,3kaxbe,2qh72,jokes,false,1441835293,https://old.reddit.com/r/Jokes/comments/3kaxbe/why_did_the_nun_get_charged_with_possession/,self.jokes,,Because she had a drug habit.,Why did the nun get charged with possession?,0
post,3kawgm,2qh72,jokes,false,1441834988,https://old.reddit.com/r/Jokes/comments/3kawgm/what_do_hurricanes_do_when_they_lose_arguments/,self.jokes,,"They storm off.

(I remembered this one when I saw the ""from when I was seven"" post)",What do hurricanes do when they lose arguments?,2
post,3katpt,2qh72,jokes,false,1441834005,https://old.reddit.com/r/Jokes/comments/3katpt/a_woman_is_at_her_fathers_deathbed/,self.jokes,,[deleted],A woman is at her father's deathbed.,1
post,3kath7,2qh72,jokes,false,1441833934,https://old.reddit.com/r/Jokes/comments/3kath7/why_do_people_like_iphone_6s_more_than_iphone_6/,self.jokes,,[deleted],Why do people like iPhone 6S more than iPhone 6?,0
post,3kasve,2qh72,jokes,false,1441833707,https://old.reddit.com/r/Jokes/comments/3kasve/ill_see_your_7_year_old_joke_and_ill_raise_you_my/,self.jokes,,Dam.,I'll see your 7 year old joke and I'll raise you my own. What did the fish say when it hit the wall?,101
post,3kasp3,2qh72,jokes,false,1441833639,https://old.reddit.com/r/Jokes/comments/3kasp3/god_i_hate_homeless_people/,self.jokes,,They make no cents... ,"God, I hate homeless people",7
post,3kasmt,2qh72,jokes,false,1441833617,https://old.reddit.com/r/Jokes/comments/3kasmt/what_do_race_car_drivers_wear_under_their_fire/,self.jokes,,Speedos !,What do race car drivers wear under their fire retardant suits?,7
post,3kascq,2qh72,jokes,false,1441833511,https://old.reddit.com/r/Jokes/comments/3kascq/a_joke_i_made_up_when_i_was_12_whats_the/,self.jokes,,"Neil Armstrong walks on the moon...

...and michael jackson fucks children. ",A joke I made up when i was 12? What's the difference between Neil Armstrong and Michael Jackson??,0
post,3kasbi,2qh72,jokes,false,1441833494,https://old.reddit.com/r/Jokes/comments/3kasbi/how_do_you_know_harry_potter_wasnt_jewish/,self.jokes,,[deleted],How do you know Harry Potter wasn't jewish?,0
post,3kar7z,2qh72,jokes,false,1441833099,https://old.reddit.com/r/Jokes/comments/3kar7z/a_woman_is_at_her_fathers_deathbed/,self.jokes,,[deleted],A woman is at her father's deathbed.,1
post,3kar5h,2qh72,jokes,false,1441833069,https://old.reddit.com/r/Jokes/comments/3kar5h/which_state_has_the_worst_asthma/,self.jokes,,Louiwheezeiana,Which state has the worst asthma?,2
post,3kaq07,2qh72,jokes,false,1441832650,https://old.reddit.com/r/Jokes/comments/3kaq07/hillary_clinton_and_donald_trump_walk_into_a_bar/,self.jokes,,"“The media is really tearing you apart for that scandal.”

Hillary: “You mean the Mexican gun running?”
Trump: “No, the other one.”

Hillary: “You mean SEAL Team 6?”
Trump: “No, the other one.”

Hillary: “You mean the State Dept. lying about Benghazi?”
Trump: “No, the other one.”

Hillary: “You mean voter fraud?”
Trump: “No, the other one.”

Hillary: “You mean the military not getting their votes counted?”
Trump: “No, the other one.”

Hillary: “The NSA monitoring our phone calls, emails and everything else?”
Trump: “No, the other one.”

Hillary: “You mean the of drones in our own country without the benefit of the law?”
Trump: “No, the other one.”

Hillary: “Giving 123 Technologies $300 Million and right after it declared bankruptcy and was sold to the Chinese?”
Trump: “No, the other one.”

Hillary: “You mean Obama arming the Muslim Brotherhood?”
Trump: “No the other one:”

Hillary: “The IRS targeting conservatives?”
Trump: “No, the other one.”

Hillary: “The DOJ spying on the press?”
Trump: “No, the other one.”

Hillary: “Sebelius shaking down health insurance executives?”
Trump: “No, the other one.”

Hillary: “Giving SOLYNDRA $500 MILLION DOLLARS and 3 months later they declared bankruptcy and then the Chinese bought it?”
Trump: “No, the other one.”

Hillary: “The NSA monitoring citizens’ phone calls, emails and everything else?”
Trump: “No, the other one.”

Hillary: “Obama’s ordering the release of nearly 10,000 illegal immigrants from jails and prisons, and falsely blaming the sequester?”
Trump: “No, the other one.”

Hillary: “Obama’s threat to impose gun control by Executive Order in order to bypass Congress?”
Trump: “No, the other one.”

Hillary: “Obama’s repeated violation of the law requiring me to submit a budget no later than the first Monday in February?”
Trump: “No, the other one.”

Hillary: “The 2012 vote where 115% of all registered voters in some counties voted 100% for Obama?”
Trump: “No, the other one.”

Hillary: “Obama’s unconstitutional recess appointments in an attempt to circumvent the Senate’s advise-and-consent role?”
Trump: “No, the other one.”

Hillary: “The State Department interfering with an Inspector General investigation on departmental sexual misconduct?”
Trump: “No, the other one.”

Hillary: “Me, The IRS, Clapper and Holder all lying to Congress?”
Trump: “No, the other one.”

Hillary: “I give up! … Oh wait, I think I got it! You mean that 65 million low-information voters who don’t pay taxes and get free stuff from taxpayers and stuck citizens again with the most pandering, corrupt administration in American history?”
Trump: “THAT’S THE ONE!”","Hillary Clinton and Donald Trump walk into a bar and grab a booth. Donald leans over, and with a smile on his face, says:",0
post,3kappy,2qh72,jokes,false,1441832548,https://old.reddit.com/r/Jokes/comments/3kappy/what_do_you_get_if_you_cross_a_joke_with_a/,self.jokes,https://www.reddit.com/r/Jokes/comments/3kappy/what_do_you_get_if_you_cross_a_joke_with_a/,,What do you get if you cross a joke with a rhetorical question?,5
post,3kapk3,2qh72,jokes,false,1441832493,https://old.reddit.com/r/Jokes/comments/3kapk3/a_man_always_comes_home_very_late_at_night_and/,self.jokes,,"and everyday he finds his wife at the door waiting for him. One time she saw a blond hair on his vest she said "" you were with a blond woman you cheater!"".So he promised her it won't happen again and got to spend the night in his house. The next day, he comes home looking like usual with a brown hair on his vest, his wife goes crazy and he manages to calm her down. Same thing next day when he comes home with a red hair on his vest. One day he came home with no hair on his vest. But his wife decided this was it! when she was asked why she said ""i'm sure he's been with a bald woman"" ",A man always comes home very late at night and drunk...,2
post,3kapcm,2qh72,jokes,false,1441832421,https://old.reddit.com/r/Jokes/comments/3kapcm/catch_up_or_catch_it/,self.jokes,,"What do you do meet an old friend?
What do you do when someone throws a ball?
What do you put on a hamburger?
What do you find in a litter box?",Catch Up or Catch It,2
post,3kap2q,2qh72,jokes,false,1441832318,https://old.reddit.com/r/Jokes/comments/3kap2q/how_did_the_hipster_burn_his_tongue/,self.jokes,,He drank the coffee before it was cool. ,How did the hipster burn his tongue?,24
post,3kaoj8,2qh72,jokes,false,1441832161,https://old.reddit.com/r/Jokes/comments/3kaoj8/whats_a_movie_where_arnold_swarzenegger_is/,self.jokes,,Preda-durrrr,What's a movie where Arnold swarzenegger is getting chased by a retarded alien?,0
post,3kao2n,2qh72,jokes,false,1441832014,https://old.reddit.com/r/Jokes/comments/3kao2n/heres_a_mind_bender_my_8_year_old_son_came_up/,self.jokes,,For camouflage.,Here's a mind bender my 8 year old son came up with: Why are trees green?,9
post,3kanb9,2qh72,jokes,false,1441831742,https://old.reddit.com/r/Jokes/comments/3kanb9/what_is_george_w_bushs_favourite_part_of_a/,self.jokes,,*Dubya Dubya Dubya*,What is George W Bush's favourite part of a website address?,0
post,3kamzr,2qh72,jokes,false,1441831630,https://old.reddit.com/r/Jokes/comments/3kamzr/how_do_you_know_you_are_at_a_gay_barbecue/,self.jokes,,The weiners taste like shit!,How do you know you are at a gay barbecue?,2
post,3kamlf,2qh72,jokes,false,1441831501,https://old.reddit.com/r/Jokes/comments/3kamlf/the_raunchy_rancher_nsfw/,self.jokes,,[deleted],The Raunchy Rancher (NSFW),1
post,3kal31,2qh72,jokes,false,1441830994,https://old.reddit.com/r/Jokes/comments/3kal31/did_you_hear_about_the_guy_who_nearly_drowned_in/,self.jokes,,He was saved by a strong currant.,Did you hear about the guy who nearly drowned in a bowl of muesli?,3
post,3kakt3,2qh72,jokes,false,1441830906,https://old.reddit.com/r/Jokes/comments/3kakt3/why_do_africans_prefer_electric_cars/,self.jokes,,Because they are mad at gas cars!,Why do Africans prefer electric cars?,0
post,3kakow,2qh72,jokes,false,1441830867,https://old.reddit.com/r/Jokes/comments/3kakow/how_do_you_bring_up_a_syrian_child/,self.jokes,,"Ram your arm down a shark's throat.

^^^Joke ^^^so ^^^dark, ^^^cops ^^^are ^^^shooting ^^^at ^^^it.",How do you bring up a Syrian child?,1
post,3kak3l,2qh72,jokes,false,1441830653,https://old.reddit.com/r/Jokes/comments/3kak3l/joke_i_heard_when_i_was_young_how_do_you_make_man/,self.jokes,,"You bake them with nuts.

(I was like 10 when I heard this joke)
",Joke I heard when I was young: How do you make man cookies?,2
post,3kajvi,2qh72,jokes,false,1441830590,https://old.reddit.com/r/Jokes/comments/3kajvi/how_is_my_penis_like_a_dead_midget/,self.jokes,,They're both a little stiff,How is my penis like a dead midget?,4
post,3kajgw,2qh72,jokes,false,1441830463,https://old.reddit.com/r/Jokes/comments/3kajgw/want_helping_coming_up_with_a_joke_that_fits_this/,self.jokes,,"[Dam Son](https://i.imgur.com/Wn3MHex.jpg)

Always sending my girlfriend corny jokes and was hoping to perfect this one with the added photo, but can't think of anything decent!",Want helping coming up with a joke that fits this.. Here's my go: What do you call an 8 year old Asian boy when he can beat Eminem in a rap battle?,0
post,3kajdp,2qh72,jokes,false,1441830432,https://old.reddit.com/r/Jokes/comments/3kajdp/what_is_8_in_plural/,self.jokes,,[deleted],What is 8 in plural?,0
post,3kaigp,2qh72,jokes,false,1441830130,https://old.reddit.com/r/Jokes/comments/3kaigp/my_little_cousin_dropped_this_one_on_me/,self.jokes,,"Me: Wow, you must've grown a foot since the last time I saw you!

Cosin: Nope, still have two!",My little cousin dropped this one on me:,10
post,3kaifs,2qh72,jokes,false,1441830121,https://old.reddit.com/r/Jokes/comments/3kaifs/have_you_heard_the_joke_about_the_man_with_no/,self.jokes,,"No? Probably a good thing, it's pretty tasteless.",Have you heard the joke about the man with no tongue?,3
post,3kahwd,2qh72,jokes,false,1441829952,https://old.reddit.com/r/Jokes/comments/3kahwd/a_flying_insect_just_flew_into_my_kitchen_and/,self.jokes,,[deleted],A flying insect just flew into my kitchen and exploded.,1
post,3kaheu,2qh72,jokes,false,1441829791,https://old.reddit.com/r/Jokes/comments/3kaheu/i_hate_dead_baby_jokes_theyre_so_old/,self.jokes,,Unlike the babies.,I hate dead baby jokes. They're so old.,0
post,3kagvi,2qh72,jokes,false,1441829609,https://old.reddit.com/r/Jokes/comments/3kagvi/what_do_you_call_a_midget_in_a_hospital_waiting/,self.jokes,,Imp-Patient!,What do you call a midget in a hospital waiting room constantly complaining about how long he's been waiting?,2
post,3kag4y,2qh72,jokes,false,1441829380,https://old.reddit.com/r/Jokes/comments/3kag4y/lahori/,self.jokes,,"Me: Where you from..??
He: From Lahore...!!
Me: Khoty k ghoshat ka taste tu bta....:D :P",#Lahori,0
post,3kafnm,2qh72,jokes,false,1441829203,https://old.reddit.com/r/Jokes/comments/3kafnm/thought_of_this_the_other_day_as_a_22_yo_how_do/,self.jokes,,You need to get ahead of lettuce,Thought of this the other day as a 22 y/o... How do you win the vegetable race?,5
post,3kaedp,2qh72,jokes,false,1441828734,https://old.reddit.com/r/Jokes/comments/3kaedp/corny_computer_jokes_why_was_the_spider_inside/,self.jokes,,He was looking for a webpage!,Corny computer jokes? Why was the spider inside the Computer?,1
post,3kaebk,2qh72,jokes,false,1441828709,https://old.reddit.com/r/Jokes/comments/3kaebk/there_was_a_soviet_clone_running_in_my_direction/,self.jokes,,He was Russian me.,There was a Soviet clone running in my direction,1
post,3kae5s,2qh72,jokes,false,1441828641,https://old.reddit.com/r/Jokes/comments/3kae5s/another_one_a_7_year_old_appreciates_why_did_the/,self.jokes,,"He was just doing his doody!

(Don't yell at me, I got it from a 7 year old)",Another one a 7 year old appreciates: Why did the anti-terrorist soldier blow up the toilet?,1
post,3kacz2,2qh72,jokes,false,1441828235,https://old.reddit.com/r/Jokes/comments/3kacz2/i_saw_a_kidnapping_today/,self.jokes,,[deleted],I saw a kidnapping today,4
post,3kacxo,2qh72,jokes,false,1441828217,https://old.reddit.com/r/Jokes/comments/3kacxo/since_were_doing_jokes_we_made_up_as_kids_heres/,self.jokes,,"Do you want to be black, or white?","Since we're doing jokes we made up as kids, here's mine: What did the World Chess Champion ask Michael Jackson?",63
post,3kacug,2qh72,jokes,false,1441828187,https://old.reddit.com/r/Jokes/comments/3kacug/a_boy_learns_some_dirty_words/,self.jokes,,"on the playground at school one day. He comes home and is shouting, ""Dick, cock, penis!"" when his mother hears him, slaps his cheek and says ""Young man, I dont ever want to hear those words come out of your mouth again."" The kid responds ""Would you rather hear them come IN my mouth?""",A boy learns some dirty words...,2
post,3kacmx,2qh72,jokes,false,1441828102,https://old.reddit.com/r/Jokes/comments/3kacmx/why_did_the_skittle_go_bowling/,self.jokes,,[deleted],Why did the skittle go bowling?,0
post,3kabqd,2qh72,jokes,false,1441827804,https://old.reddit.com/r/Jokes/comments/3kabqd/why_couldnt_the_bicycle_stand_up/,self.jokes,,Because it was two tyred..,Why couldn't the bicycle stand up?,1
post,3kabns,2qh72,jokes,false,1441827783,https://old.reddit.com/r/Jokes/comments/3kabns/i_give_you_a_joke_i_made_up_when_i_was_13/,self.jokes,,"Who's the fastest podracer in the galaxy?

Michael Chewbacca",I give you a joke I made up when I was 13,0
post,3kab7r,2qh72,jokes,false,1441827625,https://old.reddit.com/r/Jokes/comments/3kab7r/which_country_produces_the_most_fedoras/,self.jokes,,[deleted],Which country produces the most fedoras?,6
post,3kaaum,2qh72,jokes,false,1441827486,https://old.reddit.com/r/Jokes/comments/3kaaum/a_cat_walks_into_the_bar_and_asks_for_a_glass_of/,self.jokes,,"The bartender responds: '' Are you going to drink it or just knock it over on purpose?''
",A cat walks into the bar and asks for a glass of water.,0
post,3kaan4,2qh72,jokes,false,1441827408,https://old.reddit.com/r/Jokes/comments/3kaan4/whats_the_difference_between_your_mom_and_a/,self.jokes,,[deleted],whats the difference between your mom and a driveway in snowy winter?,0
post,3kaalp,2qh72,jokes,false,1441827397,https://old.reddit.com/r/Jokes/comments/3kaalp/heres_a_joke_i_just_now_made_up_at_age_40_why_did/,self.jokes,,[deleted],Here's a joke I just now made up at age 40: Why did the computer crash?,0
post,3kaaee,2qh72,jokes,false,1441827344,https://old.reddit.com/r/Jokes/comments/3kaaee/my_attempt_at_being_topical_how_do_you_know_which/,self.jokes,,[deleted],My attempt at being topical: How do you know which of your friends has the new iPhone 6s?,1
post,3kaa89,2qh72,jokes,false,1441827280,https://old.reddit.com/r/Jokes/comments/3kaa89/my_own_joke_that_im_incredibly_proud_of_what_kind/,self.jokes,,Purple Rain ,My own joke that I'm incredibly proud of: What kind of weather do Black Prince tomatoes grow best in?,2
post,3kaa2x,2qh72,jokes,false,1441827227,https://old.reddit.com/r/Jokes/comments/3kaa2x/what_is_the_easiest_way_to_kill_a_frenchman/,self.jokes,,"Break his neck by slamming down the toilet seat, while he is drinking.

- Otto von Bismarck",What is the easiest way to kill a frenchman?,1
post,3ka9ol,2qh72,jokes,false,1441827072,https://old.reddit.com/r/Jokes/comments/3ka9ol/worlds_best_joke/,self.jokes,,[deleted],World's best joke,0
post,3ka9o2,2qh72,jokes,false,1441827066,https://old.reddit.com/r/Jokes/comments/3ka9o2/what_did_the_robot_say_to_the_gas_pump/,self.jokes,,"""Take your finger out of your ear and listen to me!""

I saw this in a Highlights magazine when I was a kid.",What did the robot say to the gas pump?,1
post,3ka9f7,2qh72,jokes,false,1441826987,https://old.reddit.com/r/Jokes/comments/3ka9f7/when_was_adam_born/,self.jokes,,[deleted],When was Adam born?,0
post,3ka9ey,2qh72,jokes,false,1441826984,https://old.reddit.com/r/Jokes/comments/3ka9ey/a_man_goes_to_his_blind_doctor/,self.jokes,,"A man goes to his blind doctor to get his yearly flu vaccine.  He sits down and the receptionist calls him in to receive his vaccine.  He notices that his doctor comes walking down the hall holding a white can and tapping the wall.  He asks his doctor how he would be able to administer his vaccine and the doctor says ""I don't know. I guess it will be a shot in the dark.""",A man goes to his blind doctor.,1
post,3ka9el,2qh72,jokes,false,1441826980,https://old.reddit.com/r/Jokes/comments/3ka9el/was_helping_somebody_do_their_math_homework/,self.jokes,,"I then realized that her math teacher was a Sith Lord, because only Sith Lords deal in absolutes.",Was helping somebody do their math homework dealing with absolute values.,1
post,3ka962,2qh72,jokes,false,1441826888,https://old.reddit.com/r/Jokes/comments/3ka962/a_cat_walks_into_the_bar_and_asks_for_a_glass_of/,self.jokes,,[deleted],A cat walks into the bar and asks for a glass of water.,1
post,3ka95d,2qh72,jokes,false,1441826883,https://old.reddit.com/r/Jokes/comments/3ka95d/what_did_the_large_clock_say_to_the_small_clock/,self.jokes,,[removed],What did the large clock say to the small clock?,2
post,3ka904,2qh72,jokes,false,1441826835,https://old.reddit.com/r/Jokes/comments/3ka904/why_was_the_computer_embarrassed/,self.jokes,,"Because it has software, hardware, but no underwear!",Why was the computer embarrassed?,0
post,3ka8ip,2qh72,jokes,false,1441826686,https://old.reddit.com/r/Jokes/comments/3ka8ip/i_asked_my_father_if_hes_ever_studied_abroad/,self.jokes,,[deleted],I asked my father if he's ever studied abroad.,0
post,3ka8dw,2qh72,jokes,false,1441826636,https://old.reddit.com/r/Jokes/comments/3ka8dw/i_think_i_need_a_new_butt/,self.jokes,,...because mine has a crack in it,I think I need a new butt...,0
post,3ka8ce,2qh72,jokes,false,1441826620,https://old.reddit.com/r/Jokes/comments/3ka8ce/how_can_you_tell_which_of_your_friends_has_the/,self.jokes,,[deleted],How can you tell which of your friends has the new iPhone 6S?,0
post,3ka84o,2qh72,jokes,false,1441826541,https://old.reddit.com/r/Jokes/comments/3ka84o/my_grandma_passed_away_recently/,self.jokes,,[deleted],My grandma passed away recently..,1
post,3ka82e,2qh72,jokes,false,1441826526,https://old.reddit.com/r/Jokes/comments/3ka82e/a_cheetah_walks_slowly_out_of_the_stock_exchange/,self.jokes,,"...looking completely depressed. Two men, standing nearby having a smoke, watch the sad scene. One indicates the cheetah with his cigarette. 

""That's the third time I've seen him come out of there this week like that. Lost his retirement funds this time, I think.""

His partner shakes his head. ""A cheetah? Playing the stock exchange? What was it thinking?""

To which the other replies, ""Seriously - doesn't it know that cheetahs never prosper?""",A cheetah walks slowly out of the stock exchange...,0
post,3ka813,2qh72,jokes,false,1441826511,https://old.reddit.com/r/Jokes/comments/3ka813/what_is_the_smartest_thing_to_ever_come_out_of_a/,self.jokes,,[deleted],What is the smartest thing to ever come out of a woman's mouth?,0
post,3ka7k8,2qh72,jokes,false,1441826357,https://old.reddit.com/r/Jokes/comments/3ka7k8/what_did_the_libyan_dictators_wife_say_when_she/,self.jokes,,Muammar Gedoffame!,What did the Libyan Dictator's wife say when she didn't want to have sex?,1
post,3ka6bs,2qh72,jokes,false,1441825950,https://old.reddit.com/r/Jokes/comments/3ka6bs/what_do_you_call_two_breath_mints_that_were/,self.jokes,,Ex-pair-a-mints.,What do you call two breath mints that were turned into humans by a scientist?,1
post,3ka63m,2qh72,jokes,false,1441825876,https://old.reddit.com/r/Jokes/comments/3ka63m/i_see_your_childhood_joke_and_raise_you_mine_what/,self.jokes,,A kaleidoscope!,I see your childhood joke and raise you mine: What object crashes the most?,11
post,3ka5q3,2qh72,jokes,false,1441825743,https://old.reddit.com/r/Jokes/comments/3ka5q3/what_do_you_call_an_elephant_that_doesnt_matter/,self.jokes,,...Irrelephant.,What do you call an elephant that doesn't matter?,11
post,3ka5mw,2qh72,jokes,false,1441825709,https://old.reddit.com/r/Jokes/comments/3ka5mw/you_run_the_risk_of_getting_hearingaids_by/,self.jokes,https://www.reddit.com/r/Jokes/comments/3ka5mw/you_run_the_risk_of_getting_hearingaids_by/,,You run the risk of getting hearing-aids by sharing headphones with someone who already has them,0
post,3ka5aq,2qh72,jokes,false,1441825589,https://old.reddit.com/r/Jokes/comments/3ka5aq/two_middle_eastern_brothers_move_to_the_us/,self.jokes,,"they each make a bet over which will be more Americanized in a years time. At the end of the year the first brother says to the other ""Today I'm going to see my son play in a baseball game and after we're going to McDonalds for dinner"". The second looks at him and says ""Fuck off towel head"".",Two middle eastern brothers move to the US...,49
post,3ka4zx,2qh72,jokes,false,1441825481,https://old.reddit.com/r/Jokes/comments/3ka4zx/my_wife_said_if_this_gets_1500_upvotes/,self.jokes,,[deleted],My wife said if this gets 1500 upvotes...,0
post,3ka4qs,2qh72,jokes,false,1441825394,https://old.reddit.com/r/Jokes/comments/3ka4qs/so_a_termite_walks_into_a_bar/,self.jokes,,"...and asks, ""Hey, is the bar tender here?""",So a termite walks into a bar...,17
post,3ka4k5,2qh72,jokes,false,1441825328,https://old.reddit.com/r/Jokes/comments/3ka4k5/old_ghost_tracking_story/,self.jokes,,"So, a couple years ago, I was really into ghost tracking.  I loved the TV shows and thought I'd give it a try.  After researching the field heavily, I felt confident enough to form a task group with other investigators of the paranormal.  And so began my involvement with the Paranormal Emergency Response Team.  We became well known across town as being reliable and honest with our clients.  So much so, that after 5 years of responding to calls, we never once found an instance of actual ghosts.  I was very let down.  While the rest of the Paranormal Emergency Response Team continued working, I ended up leaving to work at a call center.  Jump ahead to a few days ago, I got a call on my private line which I had registered as being a former member of the Paranormal Emergency Response Team. The call was from some old lady who said there was something strange happening to her sink.  After work, I went over to give this lady some help.  It turned out to be a plumbing issue and there was nothing paranormal about it at all, she just wanted to ask me what her best option was.  I told her she just needed to replace one of the valves and it would be easy enough for someone to come in and fix.  Then I asked, ""why didn't you just call a plumber?""
""my son,"" she said.  ""I talked to him about the problem and he just  told me I should talk to someone with an ex-PERT opinion.""",Old Ghost Tracking Story,2
post,3ka3xu,2qh72,jokes,false,1441825087,https://old.reddit.com/r/Jokes/comments/3ka3xu/whats_the_definition_of_recursive/,self.jokes,,See recursive.,What's the definition of recursive?,3
post,3ka3ss,2qh72,jokes,false,1441825039,https://old.reddit.com/r/Jokes/comments/3ka3ss/what_did_they_call_bachs_kitchen/,self.jokes,,A feedbach system,What did they call Bach's kitchen?,1
post,3ka3rf,2qh72,jokes,false,1441825027,https://old.reddit.com/r/Jokes/comments/3ka3rf/hot_girl_in_my_apartment/,self.jokes,,"I got this hot girl back to my apartment the other day, we ripped each others clothes off and just went 
at it on the floor. 

I had her on her back and went down when she said ""David, can you take your glasses off they're digging into my thighs?""  So I took them off and we carried on. 

Minutes later she called again, ""David"" she said, ""Can you put your glasses back on please?"" 

""Why?"" I inquired.

""Because you're eating the carpet.""
",Hot girl in my apartment,8
post,3ka3ft,2qh72,jokes,false,1441824918,https://old.reddit.com/r/Jokes/comments/3ka3ft/kim_davis/,self.jokes,https://www.reddit.com/r/Jokes/comments/3ka3ft/kim_davis/,,Kim Davis,0
post,3ka3ay,2qh72,jokes,false,1441824866,https://old.reddit.com/r/Jokes/comments/3ka3ay/spanish_english_jokes_i_came_up_with_these_jokes/,self.jokes,,[deleted],Spanish English jokes... I came up with these jokes when I was learning Spanish. My friends still repeat them,0
post,3ka2s9,2qh72,jokes,false,1441824655,https://old.reddit.com/r/Jokes/comments/3ka2s9/what_do_you_call_an_unemployed_rasta/,self.jokes,,Jah Bless,What do you call an unemployed Rasta?,2
post,3ka2is,2qh72,jokes,false,1441824539,https://old.reddit.com/r/Jokes/comments/3ka2is/where_do_stoners_keep_their_money/,self.jokes,,In a joint account,Where do stoners keep their money?,6
post,3ka2hj,2qh72,jokes,false,1441824523,https://old.reddit.com/r/Jokes/comments/3ka2hj/samsung_developed_an_infinite_space_hard_drive/,self.jokes,,Only problem is they're still formatting it.,Samsung developed an infinite space hard drive.,3
post,3ka2ah,2qh72,jokes,false,1441824436,https://old.reddit.com/r/Jokes/comments/3ka2ah/what_does_the_british_monarch_do_on_the_throne/,self.jokes,,The Royal Wee.,What does the British monarch do on the throne?,2
post,3ka1y4,2qh72,jokes,false,1441824320,https://old.reddit.com/r/Jokes/comments/3ka1y4/fair_vs_unfair/,self.jokes,,If someone is fair skinned does it imply if they are darker it's unfair?,Fair Vs Unfair,1
post,3ka12d,2qh72,jokes,false,1441823974,https://old.reddit.com/r/Jokes/comments/3ka12d/i_have_a_confession_to_make_im_not_a_virgin/,self.jokes,,"A couple was on their honeymoon, lying in bed, about ready to consummate their marriage, when the new bride says to the husband, ""I have a confession to make, I'm not a virgin.""
The husband replies, ""That's no big thing in this day and age.""
The wife continues, ""Yeah, I've been with one guy.""
""Oh yeah? Who was the guy?""
""Tiger Woods.""
""Tiger Woods, the golfer?""
""Yeah.""
""Well, he's rich, famous and handsome. I can see why you went to bed with him.""
The husband and wife then make passionate love.
When they are done, the husband gets up and walks to the telephone.
""What are you doing?"" asks the wife.
The husband says, ""I'm hungry, I was going to call room service and get something to eat.""
""Tiger wouldn't do that.""
""Oh yeah? What would Tiger do?""
""He'd come back to bed and do it a second time.""
The husband puts down the phone and goes back to bed to make love a second time.
When they finish, he gets up and goes over to the phone. ""Now what are you doing?"" she asks.
The husband says, ""I'm still hungry so I was going to get room service to get something to eat.""
""Tiger wouldn't do that.""
""Oh yeah? What would Tiger do?""
""He'd come back to bed and do it again.""
The guy slams down the phone, goes back to bed, and makes love one more time.
When they finish he's tired and beat He drags himself over to the phone and starts to dial.
The wife asks, ""Are you calling room service?""
""No! I'm calling Tiger Woods. To find out what the par is for this damn hole.""","""I have a confession to make, I'm not a virgin.""",103
post,3ka0c1,2qh72,jokes,false,1441823701,https://old.reddit.com/r/Jokes/comments/3ka0c1/what_do_you_call_a_basketball_game_between_two/,self.jokes,,Juan-on-Juan,What do you call a basketball game between two Mexicans?,1
post,3ka09n,2qh72,jokes,false,1441823676,https://old.reddit.com/r/Jokes/comments/3ka09n/whats_the_difference_between_your_mom_and_the/,self.jokes,,The last time that many firefighters went down at the same time they built a memorial.,Whats the difference between your mom and the twin towers?,0
post,3ka093,2qh72,jokes,false,1441823671,https://old.reddit.com/r/Jokes/comments/3ka093/what_does_a_jihadist_say_when_he_is_taking_it/,self.jokes,,Allah mah butt,What does a jihadist say when he is taking it from behind?,0
post,3k9zw4,2qh72,jokes,false,1441823514,https://old.reddit.com/r/Jokes/comments/3k9zw4/bill_gates_meets_divine_brown/,self.jokes,,"Bill Gates meets Hugh Grant at a Hollywood party.
They are talking and Bill says, ""I've seen some great pictures of Divine Brown lately, I sure would like to get together with her!"" Hugh replies, ""Well Bill, you know ... since she gotten a little popular, her price has skyrocketed. She's charging a small fortune."" Bill said with a chuckle, ""Hugh, money's no object to me. What's her number?""

So, Hugh gives Bill her number and bill sets up a date.

They meet and after they finish, Bill is lying there in ecstasy, mumbling, ""God...now I know why you chose the name Divine.""
To which she replies, ""Thank you Bill...And now I know how you chose the name... Microsoft."" ",Bill Gates meets Divine Brown.,0
post,3k9zpr,2qh72,jokes,false,1441823447,https://old.reddit.com/r/Jokes/comments/3k9zpr/why_does_tigger_smell/,self.jokes,,"Becuase he hangs around with pooh!

Had to share my 5 year olds joke..",Why does tigger smell?,10
post,3k9zlx,2qh72,jokes,false,1441823403,https://old.reddit.com/r/Jokes/comments/3k9zlx/after_watching_todays_apple_event_i_can_confirm/,self.jokes,,"In fact, it'll be a huge 6S.","After watching today's Apple event, I can confirm the new iPhone will not be a failure.",2
post,3k9zd6,2qh72,jokes,false,1441823315,https://old.reddit.com/r/Jokes/comments/3k9zd6/mexican_firetruck/,self.jokes,,"A guy lived right on the border of Texas and Mexico. One day his house was on fire, the fire department said they were 30 minutes away. Panicking he went into Mexico and offered the fire Captain $10,000 to save his house. 

The Captain called his team, they jumped on the firetruck and went tearing across the river at 80 miles an hour, right when it looked like they were going to hit the house, the truck did a nice sideways slide coming to rest right in front of the burning house. 

After they put the fire out and saved the man's house, he asked ""What are you going to do with the money""? The Captain replied ""The first thing is to get those damn brakes fixed""!",Mexican Firetruck,1
post,3k9z1d,2qh72,jokes,false,1441823204,https://old.reddit.com/r/Jokes/comments/3k9z1d/how_does_hitler_tie_his_shoes/,self.jokes,,In little Nazis.,How does Hitler tie his shoes?,3
post,3k9yvf,2qh72,jokes,false,1441823149,https://old.reddit.com/r/Jokes/comments/3k9yvf/what_eats_everything/,self.jokes,,An Om-nomnivore,What eats everything?,3
post,3k9yqx,2qh72,jokes,false,1441823106,https://old.reddit.com/r/Jokes/comments/3k9yqx/how_do_you_tell_the_difference_between_an/,self.jokes,,[deleted],How do you tell the difference between an aligator and a crocodile?,0
post,3k9yhb,2qh72,jokes,false,1441822997,https://old.reddit.com/r/Jokes/comments/3k9yhb/my_girlfriend_is_american/,self.jokes,,I can't find her G spot but she can't find my country on a map,My girlfriend is American,0
post,3k9y5o,2qh72,jokes,false,1441822875,https://old.reddit.com/r/Jokes/comments/3k9y5o/this_just_in_famous_playboy_hugh_hefner_managed/,self.jokes,,"The police forced the friars to close down their stall, which was outside the Playboy mansion where they had been selling flowers. Said one friar, well, if it was anyone else we may have gotten away from it, but, unfortunately, only Hugh can prevent florist friars.

courtesy of Colin Mochrie",This Just In: Famous Playboy Hugh Hefner managed to successfully stop an order of monks from operating a business on his property.,1
post,3k9y07,2qh72,jokes,false,1441822831,https://old.reddit.com/r/Jokes/comments/3k9y07/how_does_a_mexican_use_liver_and_cheese_in_the/,self.jokes,,"Liver alone, cheese mine!
",How does a Mexican use 'liver' and 'cheese' in the same sentence?,1
post,3k9x1y,2qh72,jokes,false,1441822481,https://old.reddit.com/r/Jokes/comments/3k9x1y/whys_it_called_getting_an_abortion/,self.jokes,,Instead of razing your child? ,Why's it called getting an abortion...,1
post,3k9wtp,2qh72,jokes,false,1441822392,https://old.reddit.com/r/Jokes/comments/3k9wtp/what_did_the_leper_say_to_the_prostitute/,self.jokes,,Keep the tip.,What did the leper say to the prostitute?,37
post,3k9wle,2qh72,jokes,false,1441822326,https://old.reddit.com/r/Jokes/comments/3k9wle/whats_the_difference_between_my_erection_and_my/,self.jokes,,My wife actually looks forward to riding the motorcycle.,What's the difference between my erection and my motorcycle?,1
post,3k9wl1,2qh72,jokes,false,1441822323,https://old.reddit.com/r/Jokes/comments/3k9wl1/what_did_one_tectonic_plate_say_to_the_other/,self.jokes,,That was all your fault.,What did one tectonic plate say to the other after an earthquake?,2
post,3k9whl,2qh72,jokes,false,1441822287,https://old.reddit.com/r/Jokes/comments/3k9whl/how_do_you_know_when_a_women_is_pregnant/,self.jokes,,"She won't shut the fuck up about the shit she does because of the ""baby talking to her."" ",How do you know when a women is pregnant?,0
post,3k9wb2,2qh72,jokes,false,1441822216,https://old.reddit.com/r/Jokes/comments/3k9wb2/where_do_cats_go_to_meet_other_cats/,self.jokes,,A [chat](https://www.google.com/?gws_rd=ssl#q=cat+in+french) room,Where do cats go to meet other cats?,1
post,3k9way,2qh72,jokes,false,1441822215,https://old.reddit.com/r/Jokes/comments/3k9way/took_my_drivers_test_high_on_magic_mushrooms/,self.jokes,,Passed with flying colors.,Took my drivers test high on magic mushrooms.,26
post,3k9w34,2qh72,jokes,false,1441822141,https://old.reddit.com/r/Jokes/comments/3k9w34/i_met_a_rapper_the_other_day_who_told_me_he_was_a/,self.jokes,,He loved to get turnip,I met a rapper the other day who told me he was a vegetarian...,1
post,3k9w0h,2qh72,jokes,false,1441822112,https://old.reddit.com/r/Jokes/comments/3k9w0h/everyone_currently_living_on_planet_earth_is/,self.jokes,,[deleted],Everyone currently living on planet earth is attracted to me.,2
post,3k9vob,2qh72,jokes,false,1441821974,https://old.reddit.com/r/Jokes/comments/3k9vob/my_favorite_toilet_in_my_house_is_broken/,self.jokes,,Guess I'll have to make doo with my other one,My favorite toilet in my house is broken,10
post,3k9vnt,2qh72,jokes,false,1441821970,https://old.reddit.com/r/Jokes/comments/3k9vnt/what_drink_can_wrongly_convict_a_black_man/,self.jokes,,Tequila Mockingbird,What drink can wrongly convict a black man?,11
post,3k9vbb,2qh72,jokes,false,1441821844,https://old.reddit.com/r/Jokes/comments/3k9vbb/please_call_this_number/,self.jokes,,[removed],Please call this number,1
post,3k9v3x,2qh72,jokes,false,1441821781,https://old.reddit.com/r/Jokes/comments/3k9v3x/what_happened_to_the_illegally_parked_frog/,self.jokes,,It got toad away.,What happened to the illegally parked frog?,36
post,3k9uww,2qh72,jokes,false,1441821708,https://old.reddit.com/r/Jokes/comments/3k9uww/a_man_passing_through_a_rural_village_walks_into/,self.jokes,,"A man passing through a rural village walks into the local tavern. He sits down and is soon greeted by the bartender. The bartender pours him a beer as he sees the man admiring the craftsmanship of the bar.

""You see this bar?"" asks the bartender. ""I crafted this with my own two hands. I cut the timber myself, I chiseled it myself, and sanded it myself. But do you think anyone calls me Joe the Carpenter? No, no. They don't.""

The man shakes his head, sympathizing with the bartender, and continues to drink his beer as the bartender points out the window. ""You see that rock wall around the entrance?"" The man nodded. ""I built that too. I found the stone myself. I carried it all the way to town. I mixed the mortar and I laid and shaped the stone all on my own. It's a beautiful wall and I am very proud of it. But do you think anyone calls me Joe the Stonemason?"" the bartender asked, ""No! Nobody calls me that!""

""But I fuck ONE goat...""

Edit: word",A man passing through a rural village walks into the local tavern...,17
post,3k9urt,2qh72,jokes,false,1441821657,https://old.reddit.com/r/Jokes/comments/3k9urt/these_are_my_reigning_champion_twoliners/,self.jokes,,"What do you call a kingdom with a lock?

Gate Britan.

.

What do you call an opinionated island?

View Zealand.
",These are my reigning champion two-liners.,1
post,3k9uj8,2qh72,jokes,false,1441821574,https://old.reddit.com/r/Jokes/comments/3k9uj8/movies_you_wish_tom_cruise_would_star_in/,self.jokes,,Remission Impossible ,Movies you wish Tom Cruise would star in:,15
post,3k9uee,2qh72,jokes,false,1441821530,https://old.reddit.com/r/Jokes/comments/3k9uee/have_you_ever_seen_ray_chales_wife/,self.jokes,,Neither has he.,Have you ever seen Ray Chales´ Wife?,5
post,3k9txl,2qh72,jokes,false,1441821367,https://old.reddit.com/r/Jokes/comments/3k9txl/what_is_the_difference_between_a_bullet_and_a_jew/,self.jokes,,[deleted],What is the difference between a bullet and a Jew?,0
post,3k9tvx,2qh72,jokes,false,1441821348,https://old.reddit.com/r/Jokes/comments/3k9tvx/why_did_the_gay_chef_love_making_dill_crackers/,self.jokes,,Because he got to handle the dill dough.,Why did the gay chef love making dill crackers?,0
post,3k9tp6,2qh72,jokes,false,1441821290,https://old.reddit.com/r/Jokes/comments/3k9tp6/where_did_they_invent_jam/,self.jokes,,Jam maker.,Where did they invent jam?,1
post,3k9tm2,2qh72,jokes,false,1441821259,https://old.reddit.com/r/Jokes/comments/3k9tm2/i_never_use_double_negatives_irregardless_of_what/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k9tm2/i_never_use_double_negatives_irregardless_of_what/,,"I never use double negatives, irregardless of what anyone says.",0
post,3k9th0,2qh72,jokes,false,1441821209,https://old.reddit.com/r/Jokes/comments/3k9th0/why_dont_muslims_drink/,self.jokes,,Because it's not alcohalal.,Why don't Muslims drink?,2
post,3k9tf3,2qh72,jokes,false,1441821190,https://old.reddit.com/r/Jokes/comments/3k9tf3/why_cant_ray_charles_read_or_write/,self.jokes,,"Because he's dead.

If you thought this was going to be a racist or blind joke, shame on you.",Why can't Ray Charles read or write?,1
post,3k9t2a,2qh72,jokes,false,1441821048,https://old.reddit.com/r/Jokes/comments/3k9t2a/whats_the_difference_between_an_erection_and_a/,self.jokes,,I don't have a Camaro....,What's the difference between an erection and a Camaro?,2
post,3k9ssj,2qh72,jokes,false,1441820945,https://old.reddit.com/r/Jokes/comments/3k9ssj/how_to_sleep_correctly/,self.jokes,,"I have a hard time sleeping correctly so I consulted my physiotherapist on how I should be sleeping. He told me that I should be sleeping in the fetal position like when you were in the womb. But I was a C-section so I tried sleeping with a phone chord wrapped around my neck.

..Slept like a baby",How to sleep correctly?,2
post,3k9sox,2qh72,jokes,false,1441820905,https://old.reddit.com/r/Jokes/comments/3k9sox/why_did_the_shipping_company_go_under/,self.jokes,,[deleted],Why did the shipping company go under?,0
post,3k9s1n,2qh72,jokes,false,1441820682,https://old.reddit.com/r/Jokes/comments/3k9s1n/heres_a_good_one/,self.jokes,,[removed],Here's a good one.,1
post,3k9ruw,2qh72,jokes,false,1441820608,https://old.reddit.com/r/Jokes/comments/3k9ruw/james_bond_showing_his_new_watch_to_a_girl/,self.jokes,,"Bond: My watch says you are not a virgin.

Girl: But I am a virgin.

Bond: Oh my watch is 20 mins ahead.",James Bond showing his new watch to a Girl.,0
post,3k9rrv,2qh72,jokes,false,1441820575,https://old.reddit.com/r/Jokes/comments/3k9rrv/i_quit_a_job_rewriting_preclassical_greek/,self.jokes,,It feels like ancient history.,I quit a job re-writing pre-classical Greek literature into braille. This was months ago.,1
post,3k9rbp,2qh72,jokes,false,1441820415,https://old.reddit.com/r/Jokes/comments/3k9rbp/one_liner_i_made_up/,self.jokes,,I'm a depressed comedian. My life's a joke.,One liner I made up,0
post,3k9r2c,2qh72,jokes,false,1441820322,https://old.reddit.com/r/Jokes/comments/3k9r2c/waiter_waiting_for_a_tip/,self.jokes,,"A family walks into a restaurant, the waiter serves them who is exceptionally kind. He does an amazing job, treating them nicely, and even helping them with their children.

The waiter walks back into the kitchen and overhears the family saying: ""We should give him a $100 tip"" The waiter gets excited, and continues to listen. One of the family members says: ""But, I can't do it alone!"" ""Maybe we can all come together"" The family agrees.

The waiter is happy, excited, and waits anxiously for his tip. So he waits, gives the bill, and continues to wait. The family would not leave, and continued to sit at the table. An hour passed, the waiter  
could not wait anymore. So he walks up to the family.

The waiter tells them: ""Are you alright? Is there anything wrong?""
The family responds: ""When you seed $100 of evil, the roots kill 100 things around it. But when you seed $100 of good, ten thousand good prospers."" Then the family gets up, and leave. 

The man searches the table, and finds nothing, but the bill, and five dollars worth of tip.",Waiter waiting for a tip...,0
post,3k9q88,2qh72,jokes,false,1441820030,https://old.reddit.com/r/Jokes/comments/3k9q88/doctor_said_to_someone_that_smoking_is_causing/,self.jokes,, he said I am not hurry,doctor said to someone that smoking is causing slow death for you ...,1
post,3k9q4s,2qh72,jokes,false,1441819994,https://old.reddit.com/r/Jokes/comments/3k9q4s/dont_ever_buy_an_asian_computer/,self.jokes,,[deleted],Don't ever buy an Asian computer..,2
post,3k9pnm,2qh72,jokes,false,1441819819,https://old.reddit.com/r/Jokes/comments/3k9pnm/what_did_the_human_torch_tell_the_waiter_he/,self.jokes,,"Filet, mon.",What did the Human Torch tell the waiter he wanted at the Jamaican steakhouse?,1
post,3k9paj,2qh72,jokes,false,1441819692,https://old.reddit.com/r/Jokes/comments/3k9paj/the_investigation_of_ceres_was_pretty_dull_and/,self.jokes,,"Except for the discoveries in 2015, those were the two lone bright spots.",The investigation of Ceres was pretty dull and uneventful in general.,1
post,3k9nko,2qh72,jokes,false,1441819110,https://old.reddit.com/r/Jokes/comments/3k9nko/man_and_woman_on_an_airplane/,self.jokes,,"A man boarded an airplane and took his seat. As he settled in, he glanced up and saw the most beautiful woman boarding the plane. He soon realized She was heading straight towards his seat. As fate would have it, she took The seat right beside his. Eager to strike up a conversation he blurted out, “Business trip or pleasure?” She turned, smiled and said, “Business. I’m going to the Annual Nymphomaniacs of America Convention in Boston."" He swallowed hard. 

Here was the most gorgeous woman he had ever seen Sitting next to him, and she was going to a meeting of nymphomaniacs! Struggling to maintain his composure, he calmly asked, “What’s your Business at this convention?” “Lecturer,” she responded. “I use information that I have learned from my Personal experiences to debunk some of the popular myths about sexuality.” “Really?” he said. “And what kind of myths are there?” “Well,” she explained, “one popular myth is that African-American men are The most well-endowed of all men, when in fact it is the Native American Indian who is most likely to possess that trait. Another popular myth is That Frenchmen are the best lovers, when actually it is men of Mexican Descent who are the best. I have also discovered that the lover with Absolutely the best stamina is the Southern Redneck.” 

Suddenly the woman became a little uncomfortable and blushed.. “I’m Sorry,” she said, “I shouldn't really be discussing all of this with you. I don’t Even know your name.” “Tonto,” the man said, “Tonto Gonzales, but my friends call me Bubba"".",Man and woman on an airplane,18
post,3k9ngb,2qh72,jokes,false,1441819064,https://old.reddit.com/r/Jokes/comments/3k9ngb/i_can_prove_to_you_that_electronics_are_powered/,self.jokes,,by the irrefutable fact that they stop working when the smoke leaks out!,I can prove to you that electronics are powered by smoke...,5
post,3k9ndb,2qh72,jokes,false,1441819031,https://old.reddit.com/r/Jokes/comments/3k9ndb/how_soft_is_bill_gates_pillow/,self.jokes,,Microsoft.,How soft is Bill Gate's pillow?,110
post,3k9mje,2qh72,jokes,false,1441818738,https://old.reddit.com/r/Jokes/comments/3k9mje/have_you_heard_of_the_new_movie_constipation/,self.jokes,,it never came out.,Have you heard of the new movie constipation?,2
post,3k9lu9,2qh72,jokes,false,1441818499,https://old.reddit.com/r/Jokes/comments/3k9lu9/what_did_the_farmer_say_when_he_lost_his_tractor/,self.jokes,,Where's my tractor,What did the farmer say when he lost his tractor?,0
post,3k9lin,2qh72,jokes,false,1441818388,https://old.reddit.com/r/Jokes/comments/3k9lin/what_is_the_friendliest_element/,self.jokes,,Bro-mide,What is the friendliest element?,1
post,3k9ldz,2qh72,jokes,false,1441818345,https://old.reddit.com/r/Jokes/comments/3k9ldz/what_do_you_call_a_fish_with_two_knees/,self.jokes,,A tunee fish :),What do you call a fish with two knees?,3
post,3k9ldn,2qh72,jokes,false,1441818342,https://old.reddit.com/r/Jokes/comments/3k9ldn/guy_goes_to_ireland/,self.jokes,,"He is walking down a dirt path on his way to an old pub when he meets a leprechaun. He approaches the leprechaun jovially, and asks him a simple question. 
""Do rainbows always lead to a pot of gold?"" 
""Why yes they do my young sonny boy.""
""So that's why gay people are always wealthy."" ",Guy goes to Ireland,0
post,3k9l8l,2qh72,jokes,false,1441818297,https://old.reddit.com/r/Jokes/comments/3k9l8l/when_you_really_have_to_pee_and_theres_no/,self.jokes,,Urine trouble.,When you really have to pee and there's no bathroom in sight...,34
post,3k9jqb,2qh72,jokes,false,1441817763,https://old.reddit.com/r/Jokes/comments/3k9jqb/i_drive_a_delivery_truck_for_a_boss_with_an_extra/,self.jokes,,It has its UPS and downs.,I drive a delivery truck for a boss with an extra chromosome.,2
post,3k9it5,2qh72,jokes,false,1441817446,https://old.reddit.com/r/Jokes/comments/3k9it5/god_and_the_devil_were_arguing_with_each_other/,self.jokes,,"... God says to him ""I've had it! I'm taking you to court."" The devil says back ""yeah? Well where are you going to get a lawyer?"" ",God and the devil were arguing with each other...,21
post,3k9is0,2qh72,jokes,false,1441817431,https://old.reddit.com/r/Jokes/comments/3k9is0/a_pickup_like_i_thought_of_when_i_was_younger_if/,self.jokes,,On top of you. ,"A pickup like I thought of when i was younger. If I was a duck and you were a fish, and we were swimming in the same pond, what would that make me?",0
post,3k9iqd,2qh72,jokes,false,1441817409,https://old.reddit.com/r/Jokes/comments/3k9iqd/where_does_the_computer_nerd_go_for_a_drink/,self.jokes,,"At the space bar. 
How does he pay for his drinks?
Puts them on a Tab. 
Where does he do when he's had too many drinks?
The IP address. 
Where does he poop?
Install. 
How does the computer nerd potty train his son?
CTRL+P. 
",Where does the computer nerd go for a drink?,7
post,3k9iam,2qh72,jokes,false,1441817248,https://old.reddit.com/r/Jokes/comments/3k9iam/i_made_myself_golden_teeth/,self.jokes,,ro eat apples but it looks like i don't like apples,I made myself golden teeth,0
post,3k9i5l,2qh72,jokes,false,1441817200,https://old.reddit.com/r/Jokes/comments/3k9i5l/nsfwish_it_wouldve_been_my_kids_6th_birthday_today/,self.jokes,,But my pull-out game is too strong,[NSFW-ish] It would've been my kids 6th birthday today...,0
post,3k9gxk,2qh72,jokes,false,1441816772,https://old.reddit.com/r/Jokes/comments/3k9gxk/so_its_911_day_on_friday_and_i_heard_we_dont_get/,self.jokes,,[deleted],So it's 9/11 day on Friday and I heard we don't get to stay at home.,1
post,3k9g3j,2qh72,jokes,false,1441816485,https://old.reddit.com/r/Jokes/comments/3k9g3j/love_is_like_waiting_for_your_mother_to_get_off/,self.jokes,,...it never ends.,Love is like waiting for your mother to get off the phone...,4
post,3k9fft,2qh72,jokes,false,1441816235,https://old.reddit.com/r/Jokes/comments/3k9fft/the_son_of_a_farmer_start_studying_in_japan_and/,self.jokes,,[deleted],The son of a farmer start studying in Japan and send him two robots to aid in the farm,0
post,3k9fa1,2qh72,jokes,false,1441816180,https://old.reddit.com/r/Jokes/comments/3k9fa1/vote_jeb_for_president_2016/,self.jokes,,[deleted],Vote JEB for president 2016,1
post,3k9f87,2qh72,jokes,false,1441816166,https://old.reddit.com/r/Jokes/comments/3k9f87/a_trucker_who_has_been_out_on_the_road_for_two/,self.jokes,,[deleted],A trucker who has been out on the road for two weeks stops at a brothel outside Maine.,2
post,3k9f5i,2qh72,jokes,false,1441816139,https://old.reddit.com/r/Jokes/comments/3k9f5i/looking_for_a_job/,self.jokes,,[deleted],Looking for a job.,1
post,3k9e38,2qh72,jokes,false,1441815746,https://old.reddit.com/r/Jokes/comments/3k9e38/what_happened_when_the_astrophysicist_lost_a/,self.jokes,,He got a constellation prize.,What happened when the astrophysicist lost a competition?,10
post,3k9dwy,2qh72,jokes,false,1441815684,https://old.reddit.com/r/Jokes/comments/3k9dwy/i_lost_my_watch_at_a_party_once/,self.jokes,,"and then I saw a guy stepping on it while sexually harassing a girl.
I walked up to the guy and punched him right in the nose, because no one ever does that to a girl...  
Not on my watch.",I lost my watch at a party once...,448
post,3k9c5w,2qh72,jokes,false,1441815040,https://old.reddit.com/r/Jokes/comments/3k9c5w/vote_jeb_for_president_2016/,self.jokes,,Joke explain bot is always right,Vote JEB for president 2016,1
post,3k9bua,2qh72,jokes,false,1441814916,https://old.reddit.com/r/Jokes/comments/3k9bua/what_are_5_black_people_in_a_red_car/,self.jokes,,A KitKat.,What are 5 black people in a red car?,0
post,3k9ara,2qh72,jokes,false,1441814510,https://old.reddit.com/r/Jokes/comments/3k9ara/i_too_went_looking_for_secret_cove_this_morning/,self.jokes,,[deleted],I too went looking for Secret Cove this morning...,0
post,3k99ib,2qh72,jokes,false,1441814050,https://old.reddit.com/r/Jokes/comments/3k99ib/sean_connery_sylvester_stallone_and_arnold/,self.jokes,,"They are talking to the director about what roles they want to play.

Sean Connery says ""I would shertainly like to play Moshart.""

Sylvester Stallone says ""Uh, well, I guess I wanna play Beethoven.""

And so Arnold pauses a moment, and then says ""I'll be Bach.""
","Sean Connery, Sylvester Stallone, and Arnold Schwarzenegger are going to be in a movie about classical composers...",17
post,3k98sl,2qh72,jokes,false,1441813749,https://old.reddit.com/r/Jokes/comments/3k98sl/dont_ever_compete_against_heinz/,self.jokes,,You're always going to play catch up.,Don't ever compete against Heinz...,0
post,3k97t6,2qh72,jokes,false,1441813395,https://old.reddit.com/r/Jokes/comments/3k97t6/what_was_the_terrorists_pick_up_line/,self.jokes,,"'hey babe, I've got a large pipe bomb and I never pre-maturely detonate.""",What was the terrorist's pick up line?,1
post,3k97je,2qh72,jokes,false,1441813285,https://old.reddit.com/r/Jokes/comments/3k97je/today_i_have_a_test_about_irregular_verbs/,self.jokes,,[deleted],Today I have a test about irregular verbs.,1
post,3k96mv,2qh72,jokes,false,1441812945,https://old.reddit.com/r/Jokes/comments/3k96mv/eli5/,self.jokes,,Why bother... five year olds don't remember shit.  ,ELI5:,0
post,3k95jt,2qh72,jokes,false,1441812569,https://old.reddit.com/r/Jokes/comments/3k95jt/what_is_a_pedophiles_favorite_italian_meal/,self.jokes,,"Chicken Statutory....I'm going, I'm going...sorry but this is how my brain works before I've had coffee.",What is a pedophiles favorite Italian meal?,0
post,3k95e0,2qh72,jokes,false,1441812503,https://old.reddit.com/r/Jokes/comments/3k95e0/i_have_been_trying_to_lose_weight_so_ive_been/,self.jokes,,This makes it cellary.,I have been trying to lose weight so I've been keeping my junk food in the basement.,5
post,3k95d7,2qh72,jokes,false,1441812495,https://old.reddit.com/r/Jokes/comments/3k95d7/why_do_mathematician_never_go_to_the_beach/,self.jokes,,Because they got sin and cos to give them a tan,Why do mathematician never go to the beach?,11
post,3k94yw,2qh72,jokes,false,1441812355,https://old.reddit.com/r/Jokes/comments/3k94yw/what_is_michael_bays_favorite_chess_move/,self.jokes,,C4.,What is Michael Bay's favorite chess move?,20
post,3k94yc,2qh72,jokes,false,1441812348,https://old.reddit.com/r/Jokes/comments/3k94yc/johnny_shows_his_new_watch_to_his_girl_friend/,self.jokes,,"Johnny shows his new watch to his girl friend.

Johnny: My watch says you are not a virgin

Girl: But I'm still a virgin

Johnny: My watch is 20 minutes fast",Johnny shows his new watch to his girl friend,33
post,3k94ou,2qh72,jokes,false,1441812258,https://old.reddit.com/r/Jokes/comments/3k94ou/two_dust_pans_were_dry_humping/,self.jokes,,"I was like dude, get a broom already!",Two dust pans were dry humping..,5
post,3k94g1,2qh72,jokes,false,1441812164,https://old.reddit.com/r/Jokes/comments/3k94g1/what_did_the_iphone_say_to_the_fake_iphone/,self.jokes,,You're a phony,What did the iPhone say to the fake iPhone?,0
post,3k946a,2qh72,jokes,false,1441812074,https://old.reddit.com/r/Jokes/comments/3k946a/i_dont_smoke_any_more/,self.jokes,,[deleted],I don't smoke any more,1
post,3k93su,2qh72,jokes,false,1441811921,https://old.reddit.com/r/Jokes/comments/3k93su/a_computer_once_beat_me_at_chess_but_it_was_no/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k93su/a_computer_once_beat_me_at_chess_but_it_was_no/,,"A computer once beat me at chess, but it was no match for me at kick boxing. ;)",11
post,3k93p1,2qh72,jokes,false,1441811882,https://old.reddit.com/r/Jokes/comments/3k93p1/i_am_currently_working_my_ass_off_to_achieve_my/,self.jokes,, to finger my own ass while not attached to my body. ,"I am currently working my ass off to achieve my dream,",0
post,3k92xz,2qh72,jokes,false,1441811615,https://old.reddit.com/r/Jokes/comments/3k92xz/what_do_you_call_an_old_person_trying_to_fit_in/,self.jokes,,A dislocated hipster.,What do you call an old person trying to fit in with today's kids?,64
post,3k92v2,2qh72,jokes,false,1441811595,https://old.reddit.com/r/Jokes/comments/3k92v2/i_think_helen_keller_said_it_best_when_she_said/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k92v2/i_think_helen_keller_said_it_best_when_she_said/,,I think Helen Keller said it best when she said. .,0
post,3k92bg,2qh72,jokes,false,1441811379,https://old.reddit.com/r/Jokes/comments/3k92bg/husband_says_looks_like_hes_still_fucking/,self.jokes,,"Husband takes the wife to a disco. There’s a guy on the dance floor giving it large – break dancing, moon walking, back flips, the works. The wife turns to her husband and says: ""See that guy? 25 years ago he proposed to me and I turned him down."" Husband says: ""Looks like he’s still fucking celebrating!!""","Husband says: ""Looks like he’s still fucking celebrating!!""",20
post,3k92ae,2qh72,jokes,false,1441811368,https://old.reddit.com/r/Jokes/comments/3k92ae/why_is_your_nose_in_the_middle_of_your_face/,self.jokes,,It's the scenter.,Why is your nose in the middle of your face?,154
post,3k927q,2qh72,jokes,false,1441811335,https://old.reddit.com/r/Jokes/comments/3k927q/i_like_my_women_like_i_like_my_ice_cream/,self.jokes,,[deleted],"I like my women like i like my ice cream,",0
post,3k9202,2qh72,jokes,false,1441811252,https://old.reddit.com/r/Jokes/comments/3k9202/a_man_walks_into_a_psychiatrists_office_wearing/,self.jokes,,"The psychiatrist said, ""I can clearly see your nuts.""",A man walks into a psychiatrist's office wearing nothing but plastic wrap...,78
post,3k91cz,2qh72,jokes,false,1441811042,https://old.reddit.com/r/Jokes/comments/3k91cz/how_many_socialists_does_it_take_to_screw_in_a/,self.jokes,,All of them.,How many socialists does it take to screw in a lightbulb?,2
post,3k90t4,2qh72,jokes,false,1441810838,https://old.reddit.com/r/Jokes/comments/3k90t4/i_happened_to_overhear_a_guy_talking_about/,self.jokes,,"Guy 1: If I shot you in the head and you die this instant, are you sure you're gonna go to heaven?  


Guy 2: I really dont know, but Im sure you goin to hell for killing me.",I happened to overhear a guy talking about salvation to another guy...,1
post,3k90q1,2qh72,jokes,false,1441810806,https://old.reddit.com/r/Jokes/comments/3k90q1/i_dont_think_you_should_be_allowed_to_vote_if_you/,self.jokes,,[deleted],I don't think you should be allowed to vote if you don't know anything about politics. Why not?,0
post,3k909i,2qh72,jokes,false,1441810622,https://old.reddit.com/r/Jokes/comments/3k909i/car_rental_in_varanasi_new_car_rental_varanasi/,self.jokes,,[removed],Car Rental In Varanasi | New Car Rental Varanasi,1
post,3k903f,2qh72,jokes,false,1441810573,https://old.reddit.com/r/Jokes/comments/3k903f/im_going_to_make_a_movie_about_a_guy_in_a_turban/,self.jokes,,"...it'll be called ""Hyde &amp; Sikh"".",I'm going to make a movie about a guy in a turban who turns into a monster at night...,11
post,3k8zim,2qh72,jokes,false,1441810354,https://old.reddit.com/r/Jokes/comments/3k8zim/a_joke_my_philosophy_professor_told_me/,self.jokes,,"So philosophers are known to have horrible jokes, and this one is no exception. I'm just posting this for any philosophers who may or may not appreciate it. 

John has a date tomorrow with a pretty girl from his philosophy class. He's a nervous fellow and is worried about how to break the ice and start a conversation. His dad notices his son is nervous and fretting over something, and asks him what the problem is. 

""Oh dad, I have a date tomorrow and I don't know how to break the ice!"" 

""Well, son, that's easy! There are three things to talk about that will start a conversation. Food, family, and philosophy!"" 

So the next day, John goes to the ice cream parlor (it's an old joke) with his date. She stares at her ice cream and doesn't look up or speak at all. John is getting a little nervous, but remembers the ice breakers his dad taught him. 

""Do you like pizza?""

The girl looks up from her food and says ""No."" 

John, more nervous now, says ""Oh. Well do you have a brother?"" 

His date once again looks up and says ""NO!"" 

John, nervous as ever, is struggling to remember the third ice breaker his father taught him. Finally, he remembers! Philosophy! 

John straightens his face and asks ""Well, if you had a brother, would he like pizza?"" ",A joke my philosophy professor told me,69
post,3k8yre,2qh72,jokes,false,1441810059,https://old.reddit.com/r/Jokes/comments/3k8yre/an_old_lady_went_to_visit_her_dentist_when_it_was/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k8yre/an_old_lady_went_to_visit_her_dentist_when_it_was/,,"An old lady went to visit her dentist. When it was her turn, she sat in the chair, lowered her underpants, and raised her legs. The dentist said, “Excuse me, but I’m not a gynecologist.” “I know,” said the old lady. “I want you to take my husband’s teeth out.”",11
post,3k8yj0,2qh72,jokes,false,1441809971,https://old.reddit.com/r/Jokes/comments/3k8yj0/bisexuality/,self.jokes,,[deleted],Bisexuality,0
post,3k8y2e,2qh72,jokes,false,1441809785,https://old.reddit.com/r/Jokes/comments/3k8y2e/a_drunk_lady_gets_into_a_taxi/,self.jokes,,[deleted],A drunk lady gets into a taxi,1
post,3k8xt3,2qh72,jokes,false,1441809673,https://old.reddit.com/r/Jokes/comments/3k8xt3/what_did_o_say_to_q/,self.jokes,,[deleted],What did O say to Q?,5
post,3k8xnx,2qh72,jokes,false,1441809618,https://old.reddit.com/r/Jokes/comments/3k8xnx/jk_rowling_and_jk_simmons_are_getting_married/,self.jokes,,jk,JK Rowling and JK Simmons are getting married!,0
post,3k8wym,2qh72,jokes,false,1441809351,https://old.reddit.com/r/Jokes/comments/3k8wym/a_payer_for_special_needs/,self.jokes,,"

A preacher said, ""Anyone with 'special needs' who wants to be prayed over, please come forward to the front by the altar.""

With that, Leroy got in line and when it was his turn, the Preacher asked, ""Leroy, what do you want me to pray about for you?"" 

Leroy replied, ""Preacher, I need you to pray for help with my hearing."" 
The preacher put one finger of one hand in Leroy's ear, placed his other hand on top of Leroy's head and then  prayed and prayed and prayed. 
He prayed a ""blue streak"" for Leroy and the whole congregation joined in with great enthusiasm.
 
After a few minutes, the preacher removed his hands, stood back and asked, ""Leroy, how is your hearing now?""
Leroy answered, ""I don't know.  It ain't 'til next week.""

 

 

 

 

 

",A Payer for Special Needs.,62
post,3k8wy2,2qh72,jokes,false,1441809344,https://old.reddit.com/r/Jokes/comments/3k8wy2/kenny_g_walks_into_an_elevator_and_says/,self.jokes,,"“Man, this place is HAPPENING!”",Kenny G walks into an elevator and says,8
post,3k8w8f,2qh72,jokes,false,1441809063,https://old.reddit.com/r/Jokes/comments/3k8w8f/whats_the_difference_between_a_tornado_and_a/,self.jokes,,"Nothin. You're gonna lose a trailer either way.
-Robin Williams",What's the difference between a tornado and a divorce in the South?,14
post,3k8vhv,2qh72,jokes,false,1441808783,https://old.reddit.com/r/Jokes/comments/3k8vhv/why_are_blonde_jokes_always_short/,self.jokes,,So that men can understand them.,Why are blonde jokes always short?,3
post,3k8vdu,2qh72,jokes,false,1441808749,https://old.reddit.com/r/Jokes/comments/3k8vdu/i_give_to_you_a_joke_i_made_up_when_i_was_seven/,self.jokes,,"Because it had a bad driver!

*drops mic*",I give to you a joke I made up when I was seven: Why did the computer crash?,13208
post,3k8vap,2qh72,jokes,false,1441808715,https://old.reddit.com/r/Jokes/comments/3k8vap/if_you_americans_elect_donald_trump/,self.jokes,,There'll be hell toupée. ,If you Americans elect Donald Trump...,2
post,3k8v2t,2qh72,jokes,false,1441808631,https://old.reddit.com/r/Jokes/comments/3k8v2t/there_once_was/,self.jokes,,"... A man from Nebraska, 
Wait I got that part wrong, it's Alaska.
I'm awful with States,
And I'm not good with dates;
And my punch lines are just a disaster.",There once was...,2
post,3k8ury,2qh72,jokes,false,1441808524,https://old.reddit.com/r/Jokes/comments/3k8ury/why_do_celebrities_want_to_be_arctic_seaice/,self.jokes,,"Because it's getting younger, thinner and more media attention year after year.",Why do celebrities want to be Arctic sea-ice?,3
post,3k8uee,2qh72,jokes,false,1441808375,https://old.reddit.com/r/Jokes/comments/3k8uee/how_do_you_tell_if_a_redditor_was_part_of_the/,self.jokes,,[removed],How do you tell if a redditor was part of the Ellen pao lynch mob?,1
post,3k8u7k,2qh72,jokes,false,1441808305,https://old.reddit.com/r/Jokes/comments/3k8u7k/whats_the_difference_between_a_tornado_and_a/,self.jokes,,[deleted],What's the difference between a tornado and a divorce in the South?,1
post,3k8tyn,2qh72,jokes,false,1441808203,https://old.reddit.com/r/Jokes/comments/3k8tyn/a_guys_friend_has_been_on_the_toilet_for_quite_a/,self.jokes,,[deleted],A guy's friend has been on the toilet for quite a while...,1
post,3k8tjw,2qh72,jokes,false,1441808048,https://old.reddit.com/r/Jokes/comments/3k8tjw/penguins_are_scientist_by_nature/,self.jokes,,They always have to improve their slides !,Penguins are scientist by nature...,3
post,3k8scl,2qh72,jokes,false,1441807559,https://old.reddit.com/r/Jokes/comments/3k8scl/best_joke_of_all_time/,self.jokes,,[deleted],Best joke of all time.......,0
post,3k8s7y,2qh72,jokes,false,1441807505,https://old.reddit.com/r/Jokes/comments/3k8s7y/whats_the_best_holiday_to_crash_a_plain/,self.jokes,,MAY DAY! ,What's the best holiday to crash a plain?,0
post,3k8r5p,2qh72,jokes,false,1441807040,https://old.reddit.com/r/Jokes/comments/3k8r5p/have_you_ever_smelled_mothballs/,self.jokes,,How do you spread their tiny legs apart?:],Have you ever smelled mothballs?,0
post,3k8qrg,2qh72,jokes,false,1441806893,https://old.reddit.com/r/Jokes/comments/3k8qrg/whats_does_santa_clause_and_my_wife_have_in_common/,self.jokes,,They both come once every year.,What's does Santa Clause and my wife have in common?,0
post,3k8qpq,2qh72,jokes,false,1441806877,https://old.reddit.com/r/Jokes/comments/3k8qpq/bagafartcom/,self.jokes,,[removed],bagafart.com,1
post,3k8qnw,2qh72,jokes,false,1441806859,https://old.reddit.com/r/Jokes/comments/3k8qnw/an_apple_a_day_keeps_the_doctor_away/,self.jokes,, but a bowl of beans keeps everyone at bay.,"An apple a day keeps the doctor away,",2
post,3k8q9j,2qh72,jokes,false,1441806663,https://old.reddit.com/r/Jokes/comments/3k8q9j/cat_joke/,self.jokes,,"What do you call a pile of cats?



A Meowntain",Cat joke,0
post,3k8q5b,2qh72,jokes,false,1441806604,https://old.reddit.com/r/Jokes/comments/3k8q5b/a_women_is_cheating_on_her_husband_we_she_hears/,self.jokes,,"The man desperately darted around the room looking for somewhere to hide. Before he could find a good hiding space it was too late, the husband was already making his way up the staircase. Losing all hope the man hid in the bathroom. As soon as the husband arrived in the room he told his wife he going to have a shower, before she could stop him he had swung open the bathroom door, exposing the cheater. He was looking all over the room up, and down. ""Who are you?!"" asked the husband. ""Pest Control"", replied the man. ""Pest control?!"" ""for what pests?"" ""Moths"", replied the man. ""Then why are you naked?"" The naked man patted himself up and down, starred back and said ""the bastards!"" ","A women is cheating on her husband we she hears him returning. ""Quick hide!""",420
post,3k8p91,2qh72,jokes,false,1441806235,https://old.reddit.com/r/Jokes/comments/3k8p91/what_animal_is_always_ready_for_a_buffet/,self.jokes,,A platter-pus.,What animal is always ready for a buffet?,1
post,3k8np8,2qh72,jokes,false,1441805554,https://old.reddit.com/r/Jokes/comments/3k8np8/a_man_read_a_review_of_romeo_and_juliet_and_after/,self.jokes,,"Dear Mr Guyson

I'm a big fan of your magazine, and I think you have great potential as a reviewer. However, you need to put warnings for spoilers in your reviews. You've ruined Romeo and Juliet for me by giving away the ending and now I'm afraid I won't be able to see it.

Yours sincerely, John Doe.","A man read a review of Romeo and Juliet, and after getting frustrated he writes the reviewer. His letter is as follows.",0
post,3k8n67,2qh72,jokes,false,1441805310,https://old.reddit.com/r/Jokes/comments/3k8n67/i_never_let_my_kids_watch_big_band_performances/,self.jokes,,"Too much sax and violins. 




Credit to my girlfriend's dad. ",I never let my kids watch big band performances on TV.,1
post,3k8n3e,2qh72,jokes,false,1441805274,https://old.reddit.com/r/Jokes/comments/3k8n3e/i_stopped_at_a_rest_stop_to_take_a_p_now_its_a/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k8n3e/i_stopped_at_a_rest_stop_to_take_a_p_now_its_a/,,"I stopped at a rest stop to take a p, now it's a rest sto.",0
post,3k8mpt,2qh72,jokes,false,1441805093,https://old.reddit.com/r/Jokes/comments/3k8mpt/my_dr_just_diagnosed_me_as_paranoid/,self.jokes,,"Well, she didn't say that, but I know the bitch was thinking it!",My Dr. just diagnosed me as 'paranoid'!,165
post,3k8mpn,2qh72,jokes,false,1441805091,https://old.reddit.com/r/Jokes/comments/3k8mpn/there_are_three_types_of_people/,self.jokes,,People who can count and people who can't.,there are three types of people...,0
post,3k8mah,2qh72,jokes,false,1441804910,https://old.reddit.com/r/Jokes/comments/3k8mah/kim_davis_was_so_excited_to_be_released_from_jail/,self.jokes,,[deleted],Kim Davis was so excited to be released from jail.,0
post,3k8lfx,2qh72,jokes,false,1441804534,https://old.reddit.com/r/Jokes/comments/3k8lfx/iron_man_and_the_silver_surfer_should_team_up/,self.jokes,,They'd be strong alloys.,Iron Man and the Silver Surfer should team up.,63
post,3k8l48,2qh72,jokes,false,1441804376,https://old.reddit.com/r/Jokes/comments/3k8l48/she_actually_said_that/,self.jokes,,"A man was telling his buddy, ""You won't believe what happened last night... My daughter walked into the living room and said, ‘Dad, cancel my allowance immediately, forget my college tuition loan, rent my room out, throw all my clothes out the window; take my TV, and my laptop. Please take any of my jewelry to the Salvation Army or Cash Converters. Then, sell my car, take my front door key away from me and throw me out of the house. Then, disown me and never talk to me again. And don't forget to write me out of your will and leave my share to any charity you choose.’ ""

""Holy Smokes,"" replied the friend, ""she actually said that?""

""Well, she didn't put it quite like that, she actually said... 'Dad, meet my new boyfriend - Mohammed. We're going to work together on Hillary's election campaign!' ”",She actually said that?,61
post,3k8kz9,2qh72,jokes,false,1441804312,https://old.reddit.com/r/Jokes/comments/3k8kz9/whats_the_difference_between_a_virgin_and_an/,self.jokes,,[deleted],What's the difference between a virgin and an iPhone?,0
post,3k8iwg,2qh72,jokes,false,1441803386,https://old.reddit.com/r/Jokes/comments/3k8iwg/two_jungle_explorers_got_captured_by_cannibals/,self.jokes,,"Now they find themselves in a giant cauldron full of water over an open fire. The water is getting warmer and warmer and both of them realize they're done for. So they're sitting there not sure what to do when one of them lets out a chuckle. ""how could you laugh at a time like this?"" says the other one, ""we're both about to die!"".

""I know...but I just peed in their soup.""",Two jungle explorers got captured by cannibals...,106
post,3k8isa,2qh72,jokes,false,1441803341,https://old.reddit.com/r/Jokes/comments/3k8isa/this_joke_was_made_for_one_porpoise/,self.jokes,,[deleted],This joke was made for one porpoise.,0
post,3k8imh,2qh72,jokes,false,1441803265,https://old.reddit.com/r/Jokes/comments/3k8imh/a_bullet_walks_into_a_bar_depressed/,self.jokes,,"""Why the sad face?"" asks the bartender.

""I got fired.""","A bullet walks into a bar, depressed.",315
post,3k8icp,2qh72,jokes,false,1441803142,https://old.reddit.com/r/Jokes/comments/3k8icp/scotch_and_water/,self.jokes,,"A lady goes to the bar on a cruise ship and orders a scotch with two drops of water. As the bartender gives her the drink she says, ""I'm on this cruise to celebrate my 80th birthday and it's today.""

The bartender says, ""Well, since it's your birthday, I'll buy you a drink. In fact, this one is on me.""

As the woman finishes her drink the woman to her right says, ""I would like to buy you a drink, too.""

The old woman says, ""Thank you. Bartender, I want a Scotch with two drops of water.""

""Coming up,"" says the bartender.

As she finishes that drink, the man to her left says, ""I would like to buy you one, too."" The old woman says, ""Thank you. Bartender, I want another Scotch with two drops of water.""

""Coming right up,"" the bartender says.

As he gives her the drink, he says, ""Ma'am, I'm dying of curiosity. Why the Scotch with only two drops of water?""

The old woman replies, Sonny, when you're my age, you've learned how to hold your liquor... Holding your water, however, is a whole other issue.""
",Scotch and Water,16
post,3k8h42,2qh72,jokes,false,1441802588,https://old.reddit.com/r/Jokes/comments/3k8h42/why_does_the_sun_never_set_on_the_british_empire/,self.jokes,,Because God wouldn't trust an Englishman in the dark!,Why does the sun never set on the British Empire?,27
post,3k8gp9,2qh72,jokes,false,1441802396,https://old.reddit.com/r/Jokes/comments/3k8gp9/i_have_the_body_of_a_god/,self.jokes,,Buddha.,I have the body of a God.,1
post,3k8fuj,2qh72,jokes,false,1441801996,https://old.reddit.com/r/Jokes/comments/3k8fuj/why_miley_cyrus_doesnt_relate_to_hannah_montana/,self.jokes,,[deleted],Why Miley Cyrus doesn't relate to Hannah Montana anymore,0
post,3k8fd9,2qh72,jokes,false,1441801768,https://old.reddit.com/r/Jokes/comments/3k8fd9/my_best_friend_keeps_bagging_me_for_being_a_virgin/,self.jokes,,I haven't got the courage to tell him I slept with his sister.,My best friend keeps bagging me for being a virgin,3
post,3k8fc6,2qh72,jokes,false,1441801756,https://old.reddit.com/r/Jokes/comments/3k8fc6/welcome_to_jamaica_enjoy_your_stay/,self.jokes,,"A guy asks his fiance to marry him. She says okay, but only if you get a tattoo of my name on your dick. The guy agrees and gets ""Wendy"" tattooed on his dick.  When he has a soft one you could only see ""WY""

They ends up going to Jamaica for their honeymoon. The guy goes into the bathroom and sees a 7 foot Jamaican guy enters the bathroom and stands next to him taking a piss. The man looks at his dick and says ""No way, your wifes name is Wendy as well!?"". The guy looks at the man and says, ""No, it says Welcome to Jamaica enjoy your stay"".","Welcome to Jamaica, enjoy your stay",8
post,3k8faz,2qh72,jokes,false,1441801738,https://old.reddit.com/r/Jokes/comments/3k8faz/what_is_worst_then_a_repost/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k8faz/what_is_worst_then_a_repost/,,What is worst then a repost???,1
post,3k8f32,2qh72,jokes,false,1441801615,https://old.reddit.com/r/Jokes/comments/3k8f32/how_do_you_respond_when_a_jerk_rudely_brings_up_a/,self.jokes,,Douché.,How do you respond when a jerk rudely brings up a clever point?,1
post,3k8eie,2qh72,jokes,false,1441801367,https://old.reddit.com/r/Jokes/comments/3k8eie/an_intelligent_man_intelligent_woman_and_the/,self.jokes,,[deleted],"An intelligent man, intelligent woman and the tooth fairy",0
post,3k8e1k,2qh72,jokes,false,1441801124,https://old.reddit.com/r/Jokes/comments/3k8e1k/how_do_you_call_a_mexican_without_a_car/,self.jokes,,[deleted],How do you call a Mexican without a car?,0
post,3k8dav,2qh72,jokes,false,1441800793,https://old.reddit.com/r/Jokes/comments/3k8dav/last_night_i_had_a_dream_that_i_ate_a_ten_pound/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k8dav/last_night_i_had_a_dream_that_i_ate_a_ten_pound/,,"Last night I had a dream that I ate a ten pound marshmallow. When I woke up, my pillow was gone.",0
post,3k89xr,2qh72,jokes,false,1441799065,https://old.reddit.com/r/Jokes/comments/3k89xr/why_do_asian_students_do_so_well_in_school/,self.jokes,,Because an Asian without A's is a sin,Why do Asian students do so well in school?,0
post,3k89u6,2qh72,jokes,false,1441798998,https://old.reddit.com/r/Jokes/comments/3k89u6/what_did_letter_o_say_to_the_letter_q/,self.jokes,,[removed],"What did letter ""O"" say to the letter ""Q""..??",1
post,3k89jj,2qh72,jokes,false,1441798836,https://old.reddit.com/r/Jokes/comments/3k89jj/after_monday_and_tuesday_even_the_calendar_says_w/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k89jj/after_monday_and_tuesday_even_the_calendar_says_w/,,After Monday and Tuesday even the calendar says W T F.,2
post,3k89ja,2qh72,jokes,false,1441798832,https://old.reddit.com/r/Jokes/comments/3k89ja/yeh_know_these_syrians/,self.jokes,,[deleted],Yeh know these Syrians?,0
post,3k89ej,2qh72,jokes,false,1441798755,https://old.reddit.com/r/Jokes/comments/3k89ej/someone_asked_an_ex_of_dr_dre_what_did_he_do_in/,self.jokes,,"She responded, """"Beats me.""","Someone asked an ex of Dr. Dre, ""What did he do in his pastime?""",0
post,3k8934,2qh72,jokes,false,1441798587,https://old.reddit.com/r/Jokes/comments/3k8934/impact_of_movies/,self.jokes,,"Impact of Movies:

Teacher :- Who is Mahatma Gandhi?

Student:- He is the one who helped
Munna Bhai to impress his girlfriend!",Impact of Movies,0
post,3k8919,2qh72,jokes,false,1441798563,https://old.reddit.com/r/Jokes/comments/3k8919/three_men_have_to_cross_a_river_a_river_to_get/,self.jokes,,"The first man prays to God: ""Lord, oh Lord! Give me the wisdom to cross this river!"" So, God gives the man the ability to swim and he swims across. 

The second man prays to God: ""Lord, oh Lord! Give me the wisdom to cross this river!"" So, God gives the man the ability to make a raft and he crosses the river with it. 

The third man prays to God: ""Lord, oh Lord! Give me the wisdom to cross this river!"" God's getting tired by now and gives him the wisdom to cross the bridge over the river. ",Three men have to cross a river a river to get home...,1
post,3k88b8,2qh72,jokes,false,1441798155,https://old.reddit.com/r/Jokes/comments/3k88b8/what_is_never_the_answer/,self.jokes,,#,What is never the answer?,1
post,3k88aa,2qh72,jokes,false,1441798137,https://old.reddit.com/r/Jokes/comments/3k88aa/a_freudian_slip_is_when_you_say_one_thing_but/,self.jokes,,Still unsure as to whether or not that full stop adds to humorous effect.,A Freudian slip is when you say one thing but mean your mother.,26
post,3k87vd,2qh72,jokes,false,1441797896,https://old.reddit.com/r/Jokes/comments/3k87vd/why_did_u_shoot_your_wife/,self.jokes,,"Judge:why did u shoot your wife
instead of shootingher lover?

Sardar:Your honour,
it's easier to shoot a woman once,
than shooting one man every week.",Why did u shoot your wife ?,0
post,3k87lg,2qh72,jokes,false,1441797767,https://old.reddit.com/r/Jokes/comments/3k87lg/what_is_a_mexicans_favorite_queen_song/,self.jokes,," ""I Juan to break free"" ",What is a Mexican's favorite Queen song?,2
post,3k870w,2qh72,jokes,false,1441797450,https://old.reddit.com/r/Jokes/comments/3k870w/knock_knock/,self.jokes,,"You: ""Knock knock""
Victim: ""Who's there?""
You: ""I ate up""
Victim: ""I ate up who?""
(May need to be read aloud)",Knock knock,3
post,3k86cc,2qh72,jokes,false,1441797095,https://old.reddit.com/r/Jokes/comments/3k86cc/why_gordon_ramsey_hates_wwe/,self.jokes,,Because it's f*cking RAW,Why Gordon Ramsey hates WWE,36
post,3k84ml,2qh72,jokes,false,1441796105,https://old.reddit.com/r/Jokes/comments/3k84ml/i_told_my_wife_that_our_sex_tonight_will_be_out/,self.jokes,,"When she said she was sceptical, all I could say was ""I'm mixing things up, tonight my Venus is going in Uranus.""",I told my wife that our sex tonight will be out of this world.,0
post,3k823d,2qh72,jokes,false,1441794633,https://old.reddit.com/r/Jokes/comments/3k823d/i_once_told_a_girl_to_text_me_when_she_gets_home/,self.jokes,,She must have been homeless,I once told a girl to text me when she gets home,32
post,3k81ne,2qh72,jokes,false,1441794356,https://old.reddit.com/r/Jokes/comments/3k81ne/my_wife_said_all_you_do_is_talk_about_football/,self.jokes,,"There's so many more important things in life than that.

Like, what about Syria?""

I said ""Well this year I think it's between Fiorentina, Roma or Juventus",My Wife said 'All you do is talk about Football..,39
post,3k81ee,2qh72,jokes,false,1441794229,https://old.reddit.com/r/Jokes/comments/3k81ee/i_ran_into_a_fat_guy_on_the_way_to_work/,self.jokes,,Luckily I bounced back,I ran into a fat guy on the way to work,10
post,3k815y,2qh72,jokes,false,1441794099,https://old.reddit.com/r/Jokes/comments/3k815y/did_you_know_what_dr_dre_named_his_headphone/,self.jokes,,[deleted],Did you know what Dr. Dre named his headphone brand after?,0
post,3k80or,2qh72,jokes,false,1441793802,https://old.reddit.com/r/Jokes/comments/3k80or/alex_jones_is_a_joke/,self.jokes,,[removed],Alex Jones is a joke,1
post,3k7ysr,2qh72,jokes,false,1441792686,https://old.reddit.com/r/Jokes/comments/3k7ysr/how_do_you_know_when_someones_read_the_game_of/,self.jokes,,[deleted],How do you know when someone's read the Game of Thrones books?,3
post,3k7xcp,2qh72,jokes,false,1441791800,https://old.reddit.com/r/Jokes/comments/3k7xcp/how_do_you_know_when_someones_read_the_game_of/,self.jokes,,[deleted],How do you know when someone's read the Game of Thrones books?,1
post,3k7wuc,2qh72,jokes,false,1441791503,https://old.reddit.com/r/Jokes/comments/3k7wuc/whats_the_most_slippery_country/,self.jokes,,Greece.,Whats the most slippery country?,5
post,3k7ug0,2qh72,jokes,false,1441790057,https://old.reddit.com/r/Jokes/comments/3k7ug0/ama_request_kim_davis/,self.jokes,,"I would like to hear her answer this question, for she seems uniquely qualified to do so:

If a man and woman from Kentucky get a divorce, are they still brother and sister?",AMA Request: Kim Davis.,11
post,3k7uev,2qh72,jokes,false,1441790032,https://old.reddit.com/r/Jokes/comments/3k7uev/i_accidentally_dropped_my_phone_while_on_the/,self.jokes,,"Good thing it was on airplane mode, so I've got that goin' for me which is nice.  
  

Source: RyanRems",I accidentally dropped my phone while on the rooftop...,0
post,3k7te9,2qh72,jokes,false,1441789380,https://old.reddit.com/r/Jokes/comments/3k7te9/clear_before_beer_and_your_clear_to_steer/,self.jokes,,into other cars or near by pedestrians killing them and or yourself so don't fucking drink and drive you fucking moron!,"Clear before beer, and your clear to steer...",0
post,3k7tdw,2qh72,jokes,false,1441789377,https://old.reddit.com/r/Jokes/comments/3k7tdw/a_zebra_walks_into_a_bar/,self.jokes,,"He orders a drink and leaves. A few minutes later a horse walks into the bar. The bartender asks ""Hey man! What happened to your pajamas?""",A zebra walks into a bar...,1
post,3k7tbc,2qh72,jokes,false,1441789334,https://old.reddit.com/r/Jokes/comments/3k7tbc/a_14yr_old_boy_ran_into_his_house_yelling_mom_mom/,self.jokes,,"Replied the boy The mother gasped, raised her hand and slapped the boy across the face. ""get up to your room and stay ther until your father gets home!!"" yelled the mother. An hour later the boys father arrived home, got the update from the mother and went upstairs to talk to the boy. ""So I hear you had sex for the first time today"" said the father ""Your mother is upset, but I think this is something for a father and son to celebrate! What do you say we go and get you that motor-bike you've been asking for?"" ""wow, answered the boy, ""But do you think we can wait until tomorrow, my ass is still killing me!!

","A 14yr old boy ran into his house yelling ""mom mom come quick, I have great news!"" The mother asked ""what is it, what's so exciting!"" ""I had sex for the first time today!""",17
post,3k7t4a,2qh72,jokes,false,1441789185,https://old.reddit.com/r/Jokes/comments/3k7t4a/joe_was_about_to_remove_a_huge_rock_from_his_land/,self.jokes,,"-What are you doing? Thats my house. Please don't remove it, begged the gnome.
-But I would really need to move the rock.

-What if I told you that if you leave it I will grant you three wishes, but don't get to greedy, your neighbor will get twice of what you wish.

Joe really didn't like his neighbor just like you probably didn't like your worst boss.
After thinking for a while he asked the gnome.
Will it hurt a lot if I wish I only had one testicle...",Joe was about to remove a huge rock from his land when a small gnome appeared from beneath the rock.,0
post,3k7s7h,2qh72,jokes,false,1441788621,https://old.reddit.com/r/Jokes/comments/3k7s7h/why_do_people_push_the_elevator_buttons_with/,self.jokes,,[deleted],Why do people push the elevator buttons with their fingers and others with their thumbs?,0
post,3k7qon,2qh72,jokes,false,1441787707,https://old.reddit.com/r/Jokes/comments/3k7qon/how_do_you_call_a_boomerang_that_doesnt_come_back/,self.jokes,,Stick,How do you call a boomerang that doesn't come back?,1
post,3k7qd7,2qh72,jokes,false,1441787536,https://old.reddit.com/r/Jokes/comments/3k7qd7/mad_cow_disease_jokes/,self.jokes,,"So there were these two cows, chatting over the fence
between their fields.
The first cow said,""I tell you, this mad-cow-disease is really
pretty scary. They say it is spreading fast; I heard it hit
some cows down on the Johnson Farm.""
The other cow replies, ""Hell, I ain't worried, it don't affect us
ducks.""
A female reporter was conducting an interview with a farmer
about Mad Cow Disease. ""Mr. Brown, do you have any idea
what might be the cause of the disease?""
""Sure. Do you know the bulls only screw the cows once a
year?""
""Umm, sir, that is a new piece of information, but what's the
relationship between this and Mad Cow?""
""And did you know we milk the cows twice a day?""
""Mr. Brown, that's interesting, but, what's the point?""
""Lady, the point is this: if I'm playing with your tits twice a
day, but only screwing you once a year, wouldn't you go
mad, too?""
",Mad cow disease jokes,0
post,3k7q8f,2qh72,jokes,false,1441787454,https://old.reddit.com/r/Jokes/comments/3k7q8f/new_channels_bin_laden_dead/,self.jokes,," That's ruined the game, what do we do now it's our turn to hide? ",New Channels: Bin Laden dead,0
post,3k7pib,2qh72,jokes,false,1441787002,https://old.reddit.com/r/Jokes/comments/3k7pib/since_were_at_it_dating_in_your_30s_is_like/,self.jokes,,The good ones are all taken. But you can always get one from an exotic country...,Since we're at it: Dating in your 30s is like registering a domain name...,16
post,3k7p53,2qh72,jokes,false,1441786761,https://old.reddit.com/r/Jokes/comments/3k7p53/what_do_you_call_it_when_a_banana_eats_another/,self.jokes,,Canabananalism,What do you call it when a banana eats another banana?,10
post,3k7oy7,2qh72,jokes,false,1441786642,https://old.reddit.com/r/Jokes/comments/3k7oy7/what_happened_to_the_two_gladiator_olives/,self.jokes,,They were pitted against each other,What happened to the two gladiator olives?,3
post,3k7myq,2qh72,jokes,false,1441785417,https://old.reddit.com/r/Jokes/comments/3k7myq/so_i_saw_a_boy_at_the_shops_today_on_his_own/,self.jokes,,"It looked like fun and he seemed lonely so I joined in with him. 
Nek minnit his parents come over spitting chips!
Turns out he has cerebral palsy and I'm a terrible person.","So I saw a boy at the shops today on his own, pretending to be a dinosaur.",0
post,3k7m7q,2qh72,jokes,false,1441784977,https://old.reddit.com/r/Jokes/comments/3k7m7q/what_is_it_called_when_you_kill_a_friend/,self.jokes,,Homiecide.... I'll^see^myself^out...,What is it called when you kill a friend?,3
post,3k7jd4,2qh72,jokes,false,1441783360,https://old.reddit.com/r/Jokes/comments/3k7jd4/i_was_making_a_graph_of_my_past_relationships/,self.jokes,,Full disclosure: I saw this in yik yak thought is share it here. :) ,I was making a graph of my past relationships. First I drew the Ex axis then the Why axis.,4
post,3k7isl,2qh72,jokes,false,1441783007,https://old.reddit.com/r/Jokes/comments/3k7isl/whats_the_definition_of_a_will/,self.jokes,,"(Come on, it's a dead giveaway!)",What's the definition of a will?,21
post,3k7hoj,2qh72,jokes,false,1441782385,https://old.reddit.com/r/Jokes/comments/3k7hoj/i_asked_the_waitress_if_she_wanted_a_good_tip_and/,self.jokes,,She said: Just the tip.,I asked the waitress if she wanted a good tip and a quickie.,4
post,3k7hcw,2qh72,jokes,false,1441782201,https://old.reddit.com/r/Jokes/comments/3k7hcw/my_wife_cant_cook_so_she_asked_me_for_help_in/,self.jokes,,She put one in the bedroom and one in the bathroom.. Ijit.,My wife can't cook so she asked me for help in baking a cake. I told her to separate 2 eggs...,2
post,3k7gf8,2qh72,jokes,false,1441781672,https://old.reddit.com/r/Jokes/comments/3k7gf8/im_not_saying_i_have_a_small_dick/,self.jokes,,[deleted],I'm not saying I have a small dick,0
post,3k7f55,2qh72,jokes,false,1441780906,https://old.reddit.com/r/Jokes/comments/3k7f55/two_men_walk_into_a_bar/,self.jokes,,Well that wasn't very smart,Two men walk into a bar,0
post,3k7dkt,2qh72,jokes,false,1441780098,https://old.reddit.com/r/Jokes/comments/3k7dkt/been_reading_about_instinctive_behaviors/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k7dkt/been_reading_about_instinctive_behaviors/,,"Been reading about instinctive behaviors. Apparently, my natural reaction to seeing an attractive woman is a Fixed Action Pattern (in short, FAP).",7
post,3k7ary,2qh72,jokes,false,1441778608,https://old.reddit.com/r/Jokes/comments/3k7ary/whats_6_inches_long_2_inches_wide_and_drives/,self.jokes,,[deleted],"What's 6 inches long, 2 inches wide and drives women wild?",0
post,3k7a20,2qh72,jokes,false,1441778240,https://old.reddit.com/r/Jokes/comments/3k7a20/theres_only_one_thing_i_love_more_than_bacon/,self.jokes,,...and I can't put pussy in my mashed potatoes. ,There's only one thing I love more than bacon,6
post,3k79yp,2qh72,jokes,false,1441778195,https://old.reddit.com/r/Jokes/comments/3k79yp/my_bumper_sticker_says_honk_if_you_think_im_sexy/,self.jokes,,[deleted],"My bumper sticker says ""Honk if you think I'm sexy""",430
post,3k79ox,2qh72,jokes,false,1441778056,https://old.reddit.com/r/Jokes/comments/3k79ox/i_wasnt_sure_about_my_beard_at_first/,self.jokes,,[deleted],I wasn't sure about my beard at first...,0
post,3k7975,2qh72,jokes,false,1441777780,https://old.reddit.com/r/Jokes/comments/3k7975/a_black_woman_had_5_sons_name_tyrone_tyrone/,self.jokes,,"How did she tell them apart?


She called them by their last names","A black woman had 5 sons name Tyrone, Tyrone, Tyrone, Tyrone and Tyrone....",60
post,3k78y9,2qh72,jokes,false,1441777627,https://old.reddit.com/r/Jokes/comments/3k78y9/what_is_brown_and_rhymes_with_snoop_dogg/,self.jokes,,Dr. Dre,What is brown and rhymes with snoop dogg?,3
post,3k78ay,2qh72,jokes,false,1441777271,https://old.reddit.com/r/Jokes/comments/3k78ay/a_redditor_sees_a_comment_that_he_doesnt_agree/,self.jokes,,...and gives it an upvote because it's a valid point. ,A Redditor sees a comment that he doesn't agree with...,71
post,3k77a3,2qh72,jokes,false,1441776689,https://old.reddit.com/r/Jokes/comments/3k77a3/what_is_the_difference_between_a_black_man_and_an/,self.jokes,,An elevator can raise a child.,What is the difference between a black man and an elevator?,0
post,3k768b,2qh72,jokes,false,1441776155,https://old.reddit.com/r/Jokes/comments/3k768b/these_daysbots_like_siri_pretend_to_be_human/,self.jokes,,[deleted],"These days,bots, like Siri, pretend to be human beings, and human beings...",0
post,3k73o9,2qh72,jokes,false,1441774896,https://old.reddit.com/r/Jokes/comments/3k73o9/cs_go_joke/,self.jokes,,"How many CS GO silver ranked players does it take to fix a light bulb.

None cause they cant climb the ladder ahahahahahaha ",Cs go joke,6
post,3k739s,2qh72,jokes,false,1441774722,https://old.reddit.com/r/Jokes/comments/3k739s/whats_helen_kellers_favorite_color/,self.jokes,,[deleted],What's Helen Keller's favorite color?,2
post,3k72i1,2qh72,jokes,false,1441774327,https://old.reddit.com/r/Jokes/comments/3k72i1/what_are_rich_people_called_in_japan/,self.jokes,,Milyennaires,What are rich people called in Japan?,0
post,3k72dw,2qh72,jokes,false,1441774263,https://old.reddit.com/r/Jokes/comments/3k72dw/whats_the_definition_of_a_will/,self.jokes,,[deleted],What's the definition of a will?,0
post,3k71zg,2qh72,jokes,false,1441774103,https://old.reddit.com/r/Jokes/comments/3k71zg/2_mexican_brothers_crossed_the_border_and_need/,self.jokes,,"(Slightly Racist - You have been warned)

Jose and Juan, 2 brothers, crossed the border to USA and had no cash. Their plan was to beg on the streets for some money. So the two brothers both got cardboard and made their own signs. Juan says ""Lets split up, you go up the street, I do down, we meet here at night.""

Jose agrees to the plan and heads up the street with his sign begging for money at a busy intersection. Juan feeling good about his plan goes down the street at another intersection and begs also.

By the end of the day, the 2 brothers meet where they started with all their money. Juan, still feeling good about his plan, shows his younger brother he made $40! While Juan is laughing, his younger brother pulls out $200 from his pockets. 

Juan shocked ask his brother, ""How did you make so much money?"" His brother responded, ""Read my sign."" Jose's sign reads ""Need $20 to go back to Mexico""

(My dad told me this joke when I was 10, I live in LA area)",2 Mexican brothers crossed the border and need money,118
post,3k71vf,2qh72,jokes,false,1441774042,https://old.reddit.com/r/Jokes/comments/3k71vf/why_did_the_otter_cross_the_road/,self.jokes,,To get to the OTTER side!,Why did the otter cross the road?,0
post,3k70lm,2qh72,jokes,false,1441773486,https://old.reddit.com/r/Jokes/comments/3k70lm/your_greatest_puns/,self.jokes,,"Please, I love puns. Lots of puns. Any kind. Bring em on!",Your greatest puns!,0
post,3k70ep,2qh72,jokes,false,1441773395,https://old.reddit.com/r/Jokes/comments/3k70ep/why_does_isis_wear_condoms_when_they_have_sex/,self.jokes,,So they can fuck two goats at once! ,Why does ISIS wear condoms when they have sex?,0
post,3k6zn4,2qh72,jokes,false,1441773050,https://old.reddit.com/r/Jokes/comments/3k6zn4/whats_the_difference_between_a_catfish_and_a/,self.jokes,,"One is a filthy, slimy, bottom-feeding, scum-sucking monstrosity with long whiskers, and the other is a fish.",What's the difference between a catfish and a Frenchman?,2
post,3k6zm3,2qh72,jokes,false,1441773033,https://old.reddit.com/r/Jokes/comments/3k6zm3/my_girlfriend_told_me_to_go_out_and_bring_back/,self.jokes,,I came home drunk.,My girlfriend told me to go out and bring back something that made her look sexy.,11
post,3k6zak,2qh72,jokes,false,1441772864,https://old.reddit.com/r/Jokes/comments/3k6zak/tell_me_something_a_farmer_cares_more_about_than/,self.jokes,,[deleted],Tell me something a farmer cares more about than his wife?,3
post,3k6yoy,2qh72,jokes,false,1441772599,https://old.reddit.com/r/Jokes/comments/3k6yoy/my_girlfriend_treats_me_like_a_god/,self.jokes,,She ignores me until she needs something.,My girlfriend treats me like a god.,7
post,3k6yai,2qh72,jokes,false,1441772409,https://old.reddit.com/r/Jokes/comments/3k6yai/an_englishman_a_frenchman_and_joseph_stalin_are/,self.jokes,,"and they spot a beautiful portrait of Adam and Eve.

""Oh, look how dignified and noble they are! It's clear that Adam and Eve were English"", says the Englishman.

""No way, man! Observe their grace and beauty and love! They are clearly French!"", says the Frenchman.

The two keep arguing until Stalin simply scoffs and laughs while shaking his head. ""Comrades, you are missing the point! Look at them. They have no clothes and no shelter, and they have only apples to eat, yet they are told that they are living in paradise. They are obviously Russian!"".","An Englishman, a Frenchman, and Joseph Stalin are in an art exhibit",14
post,3k6xd2,2qh72,jokes,false,1441772014,https://old.reddit.com/r/Jokes/comments/3k6xd2/what_do_you_get_when_you_cross_pewdiepie_and/,self.jokes,,[deleted],What do you get when you cross pewdiepie and youtube?,0
post,3k6xam,2qh72,jokes,false,1441771982,https://old.reddit.com/r/Jokes/comments/3k6xam/id_also_tell_you_a_joke_about_how_my_balls_hang/,self.jokes,,But that's too low.,I'd also tell you a joke about how my balls hang. . .,0
post,3k6x1z,2qh72,jokes,false,1441771861,https://old.reddit.com/r/Jokes/comments/3k6x1z/how_many_trolls_does_it_take_to_read_a_joke/,self.jokes,,None.  They get chumps like you to do it.  CHUMPS.,How many trolls does it take to read a joke.,0
post,3k6wuc,2qh72,jokes,false,1441771759,https://old.reddit.com/r/Jokes/comments/3k6wuc/hillary_clinton_the_pope_barack_obama_and_a_boy/,self.jokes,,"and the plane is crashing!

There are three parachutes that the four can use, but each parachute can only carry one person.

""As the leader of the free world, I'm afraid I must insist that I take a parachute. All of America depends on me!"", says Barack Obama, and he is given a parachute.

After he jumps, Hillary Clinton goes next. ""I am the most gifted and most intelligent woman in all of creation and I am America's future president, so I DEMAND a parachute!"". The boy sighs and hands her it, and she jumps out of the window.

Finally, only the Pope and the boy scout are left.

""My child, I have already lived a long and gifted life, and I am ready to join the Lord in Heaven, so take the parachute."", the Pope says.

""You take one."", says the boy.

""No, you do not understand. I am not long for this earth anyway and am ready to sacrifice my elderly self for you so you can live out your life."", says the Pope.

""No, really, you take a parachute!"", says the boy scout.

""Son, we don't have much time! There is only one parachute left and you must take it."", says the Pope.

""No, we have two parachutes! I gave that bitch my backpack!""","Hillary Clinton, the Pope, Barack Obama, and a boy scout are all on a plane",84
post,3k6wb4,2qh72,jokes,false,1441771534,https://old.reddit.com/r/Jokes/comments/3k6wb4/why_would_you_throw_a_rock_at_a_mexican_man/,self.jokes,,"Because it's probably your bike. 

Why would you throw a rock at a black man riding a bike? 

Because it's probably your black man.",Why would you throw a rock at a Mexican man riding a bike?,0
post,3k6vtx,2qh72,jokes,false,1441771291,https://old.reddit.com/r/Jokes/comments/3k6vtx/i_prefer_oneliners/,self.jokes,,[deleted],I prefer one-liners..,0
post,3k6vom,2qh72,jokes,false,1441771218,https://old.reddit.com/r/Jokes/comments/3k6vom/id_tell_you_a_joke_about_my_penis/,self.jokes,,But it's too short &amp; not many people get it.,I'd tell you a joke about my penis. . .,2
post,3k6vlh,2qh72,jokes,false,1441771181,https://old.reddit.com/r/Jokes/comments/3k6vlh/whats_it_called_when_you_go_around_looking_for/,self.jokes,,Antiquing.,What's it called when you go around looking for stuff to buy that's made in America?,13
post,3k6vhb,2qh72,jokes,false,1441771152,https://old.reddit.com/r/Jokes/comments/3k6vhb/so_the_french_army_has_recently_installed/,self.jokes,,"That way, they can watch the fighting!",So the French army has recently installed rearview mirrors to their tanks.,34
post,3k6ty3,2qh72,jokes,false,1441770489,https://old.reddit.com/r/Jokes/comments/3k6ty3/_/,self.jokes,,[removed],:),1
post,3k6te2,2qh72,jokes,false,1441770262,https://old.reddit.com/r/Jokes/comments/3k6te2/if_i_eat_lots_of_preservatives_wont_i_live_longer/,self.jokes,,"No, but you will have a longer shelf life.
","If I eat lots of preservatives, won't I live longer?",1
post,3k6t5e,2qh72,jokes,false,1441770148,https://old.reddit.com/r/Jokes/comments/3k6t5e/what_do_you_call_a_nautical_plunderer_who_assists/,self.jokes,,A co-pirate,What do you call a nautical plunderer who assists with the flight of an aircraft?,7
post,3k6t53,2qh72,jokes,false,1441770143,https://old.reddit.com/r/Jokes/comments/3k6t53/why_do_mules_not_work_as_hard_as_horses/,self.jokes,,Because they're half-assed!,Why do mules not work as hard as horses?,1
post,3k6sea,2qh72,jokes,false,1441769872,https://old.reddit.com/r/Jokes/comments/3k6sea/some_people_say_i_have_no_soul/,self.jokes,,[deleted],Some people say I have no soul.,0
post,3k6rpv,2qh72,jokes,false,1441769606,https://old.reddit.com/r/Jokes/comments/3k6rpv/microsoft_tech_support_called_me_last_night/,self.jokes,,"as a indian, I said ""Sorry your calling Indian Tech Support""",Microsoft tech support called me last night,0
post,3k6r5c,2qh72,jokes,false,1441769385,https://old.reddit.com/r/Jokes/comments/3k6r5c/not_exactly_a_joke_but_a_funny_retort_of_my/,self.jokes,,[deleted],Not exactly a joke but a funny retort of my brothers.,1
post,3k6r3g,2qh72,jokes,false,1441769368,https://old.reddit.com/r/Jokes/comments/3k6r3g/lpt_do_not_fall_in_love_with_tennis_players/,self.jokes,,Love means nothing to them,LPT: Do not fall in love with tennis players,3
post,3k6qzq,2qh72,jokes,false,1441769324,https://old.reddit.com/r/Jokes/comments/3k6qzq/a_zoologist_a_statistician_and_a_mathematician/,self.jokes,,"While they are sitting there they see two people enter the house. A short while later they see three people leave the house.

The zoologist says ""They must have reproduced.""
The statistician says ""Our initial count must have been wrong.""
The mathematician says ""If one more person goes into that house it will be empty again.""","A zoologist, a statistician, and a mathematician are sitting across the street from an empty house.",27
post,3k6px7,2qh72,jokes,false,1441768915,https://old.reddit.com/r/Jokes/comments/3k6px7/why_did_the_chicken_cross_the_road/,self.jokes,,So I can have an opportunity to make small talk,Why did the chicken cross the road?,3
post,3k6ptw,2qh72,jokes,false,1441768879,https://old.reddit.com/r/Jokes/comments/3k6ptw/im_going_to_heaven/,self.jokes,,"Gay sex prevents abortions, suck dick for Jesus !!",I'm going to heaven,0
post,3k6pqt,2qh72,jokes,false,1441768847,https://old.reddit.com/r/Jokes/comments/3k6pqt/a_rich_man_and_a_poor_man_have_the_same_wedding/,self.jokes,,"They're both at Madison Avenue shopping for their wives. Poor man says to the Rich man, ""What'd you get your wife this year?""

He says, ""A Mercedes and a huge diamond ring."" The poor man says, ""Why'd you get her both?"" The Rich man says, ""If she doesn't like the ring, she can take it back to store in her new car, come home and still be happy."" The Poor man says, ""O.K. That works.""

The Rich man says, ""Well what did you get your wife?"" The Poor man says, ""A pair of slippers and a dildo.""

The Rich man says, ""Why'd you get her a pair of slippers and a dildo?""

The Poor man says, ""If she doesn't like the slippers, she can go fuck herself!""

Source: Tony Soprano",A rich man and a poor man have the same wedding anniversary.,3
post,3k6p3d,2qh72,jokes,false,1441768585,https://old.reddit.com/r/Jokes/comments/3k6p3d/how_do_you_know_if_your_wine_was_made_in_the_90s/,self.jokes,,It smells like teen spirit.,How do you know if your wine was made in the 90's?,1
post,3k6osl,2qh72,jokes,false,1441768469,https://old.reddit.com/r/Jokes/comments/3k6osl/wanna_hear_a_joke_about_pizza/,self.jokes,,"never mind, it's too cheesy. 

















-__-",Wanna hear a joke about pizza?,5
post,3k6oo1,2qh72,jokes,false,1441768432,https://old.reddit.com/r/Jokes/comments/3k6oo1/what_do_you_call_a_midget_fortune_teller_running/,self.jokes,,A small medium at large.,What do you call a midget fortune teller running from the police?,0
post,3k6mw9,2qh72,jokes,false,1441767689,https://old.reddit.com/r/Jokes/comments/3k6mw9/what_do_you_call_fast_food_emergencies/,self.jokes,,"Emergen-cheese.

:3",What do you call fast food emergencies?,0
post,3k6mdi,2qh72,jokes,false,1441767478,https://old.reddit.com/r/Jokes/comments/3k6mdi/what_kind_of_currency_do_aliens_use/,self.jokes,,[deleted],What kind of currency do aliens use?,0
post,3k6lno,2qh72,jokes,false,1441767196,https://old.reddit.com/r/Jokes/comments/3k6lno/what_did_michael_jackson_say_to_the_catholic/,self.jokes,,[deleted],What did Michael Jackson say to the Catholic priest?,0
post,3k6lcf,2qh72,jokes,false,1441767045,https://old.reddit.com/r/Jokes/comments/3k6lcf/a_scoliosis_patient_had_given_up_hope_of_recovery/,self.jokes,,"But after the long and painful surgery, he took his first steps and humbly said ""I stand corrected"".",A scoliosis patient had given up hope of recovery..,19
post,3k6l01,2qh72,jokes,false,1441766904,https://old.reddit.com/r/Jokes/comments/3k6l01/so_an_openly_gay_guy_patronized_a_store_in_indiana/,self.jokes,,.,So an openly gay guy patronized a store in Indiana,0
post,3k6kek,2qh72,jokes,false,1441766682,https://old.reddit.com/r/Jokes/comments/3k6kek/what_do_you_call_a_sleepwalking_nun/,self.jokes,,A roamin' Catholic.,What do you call a sleepwalking nun?,1
post,3k6hu8,2qh72,jokes,false,1441765684,https://old.reddit.com/r/Jokes/comments/3k6hu8/did_you_hear_about/,self.jokes,,"The dad who put gasoline in his daughter's sippy cup?

Doctor's say she's going to be fine. She just had a little gas.",Did you hear about...?,0
post,3k6hoc,2qh72,jokes,false,1441765618,https://old.reddit.com/r/Jokes/comments/3k6hoc/no_matter_how_bad_your_mood_is_no_matter_how_fd/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k6hoc/no_matter_how_bad_your_mood_is_no_matter_how_fd/,,"No matter how bad your mood is, no matter how f****d up you're in your life, there are still some people. Yeah ""some people"". Who can unknowingly bring that smile back on your face just by their words.",0
post,3k6fqh,2qh72,jokes,false,1441764856,https://old.reddit.com/r/Jokes/comments/3k6fqh/test_boast_please_ignore/,self.jokes,,I just hacked my friend's reddit account.,"Test boast, please ignore.",0
post,3k6fq5,2qh72,jokes,false,1441764851,https://old.reddit.com/r/Jokes/comments/3k6fq5/mayweatherfloyd_mayweather_jr_vs_andre_berto/,self.jokes,,[removed],[[Mayweather]]Floyd Mayweather Jr vs. Andre Berto Stream..Live.,1
post,3k6fl2,2qh72,jokes,false,1441764793,https://old.reddit.com/r/Jokes/comments/3k6fl2/what_do_you_think_about_euthanasia/,self.jokes,,[deleted],What do you think about euthanasia?,1
post,3k6fbb,2qh72,jokes,false,1441764675,https://old.reddit.com/r/Jokes/comments/3k6fbb/what_do_you_call_a_crocodile_who_always_lies/,self.jokes,,A croc o' shit.,What do you call a crocodile who always lies?,7
post,3k6f5e,2qh72,jokes,false,1441764605,https://old.reddit.com/r/Jokes/comments/3k6f5e/did_you_hear_about_the_epileptic_midget_who_works/,self.jokes,,They call him Little Seizures.  ,Did you hear about the epileptic midget who works at the pizzeria?,49
post,3k6eux,2qh72,jokes,false,1441764487,https://old.reddit.com/r/Jokes/comments/3k6eux/an_extremely_close_friend_just_confided_in_me/,self.jokes,,He is no longer my close friend.,An extremely close friend just confided in me that he likes comic sans.,0
post,3k6ekn,2qh72,jokes,false,1441764378,https://old.reddit.com/r/Jokes/comments/3k6ekn/i_was_opposed_when_my_wife_brought_up_the_idea_of/,self.jokes,,But my hands were tied.,I was opposed when my wife brought up the idea of trying BDSM...,1
post,3k6dm0,2qh72,jokes,false,1441763964,https://old.reddit.com/r/Jokes/comments/3k6dm0/what_is_the_difference_between_an_engineer/,self.jokes,,"An engineer is someone who comes up with equations that model reality.

A physicist is someone who comes up with a reality that models their equations.

A mathematician doesn't care.","What is the difference between an engineer, physicist, and a mathematician?",0
post,3k6d5p,2qh72,jokes,false,1441763804,https://old.reddit.com/r/Jokes/comments/3k6d5p/what_do_you_get_when_you_cross_a_joke_with_a/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k6d5p/what_do_you_get_when_you_cross_a_joke_with_a/,,What do you get when you cross a joke with a rhetorical question?,30
post,3k6csf,2qh72,jokes,false,1441763645,https://old.reddit.com/r/Jokes/comments/3k6csf/why_doesnt_barbie_have_a_family/,self.jokes,,Because Ken comes in another box. ,Why doesn't Barbie have a family?,4
post,3k6cik,2qh72,jokes,false,1441763524,https://old.reddit.com/r/Jokes/comments/3k6cik/a_man_walks_into_a_brothel_but_doesnt_have_much/,self.jokes,,[deleted],"A man walks into a brothel, but doesn't have much money",0
post,3k6blq,2qh72,jokes,false,1441763179,https://old.reddit.com/r/Jokes/comments/3k6blq/three_men_go_to_heaven_and_st_peter_says_they_are/,self.jokes,,"...so they are transported down to hell. The devil, being a reasonable guy, apologizes for the mistake, and promises to set each man up with a room filled with whatever they want. The first man asks for a room full of chocolate, which the devil procures, and closes the door behind him. The second man asks for a room full of beautiful women, the devil agrees, and shows him into the room. The third man requests a room full of Marijuana. The devil shows him in, and says ""Ok, I'll check on you in 10,000 years.""

When the devil comes back, he open the first day to find a huge fat man, covered in chocolate, and enjoying himself. He open the second door, and sees a bunch of pregnant women, and babies. 

When the devil open the third door, the man jumps out, and grabs the devil by the collar. He screams: 

""GOT A LIGHT?""","Three men go to heaven, and St. Peter says they are full....",61
post,3k6bja,2qh72,jokes,false,1441763155,https://old.reddit.com/r/Jokes/comments/3k6bja/whats_an_arborists_favorite_side_dish/,self.jokes,,Can o' peas.,What's an arborists favorite side dish?,0
post,3k6bb8,2qh72,jokes,false,1441763055,https://old.reddit.com/r/Jokes/comments/3k6bb8/my_drug_dealer_is_so_funny/,self.jokes,,[removed],my drug dealer is so funny,1
post,3k6b62,2qh72,jokes,false,1441762994,https://old.reddit.com/r/Jokes/comments/3k6b62/ironic/,self.jokes,,"One bright day in the middle of the night
Two dead boys got up to fight.
Back to back they faced each other 
Drew their swords and shot each other. 
A deaf policeman heard the noise 
and ran to save the two dead boys.
And if you don't believe it's true 
go ask the blind man, he saw it too.",Ironic,6
post,3k6ay4,2qh72,jokes,false,1441762908,https://old.reddit.com/r/Jokes/comments/3k6ay4/a_man_walked_into_a_brothel_but_doesnt_have_much/,self.jokes,,[deleted],"A man walked into a brothel, but doesn't have much money to spend",1
post,3k6an5,2qh72,jokes,false,1441762780,https://old.reddit.com/r/Jokes/comments/3k6an5/when_tim_tebow_found_out_he_got_cut_by_the_eagles/,self.jokes,,.. And even that got intercepted. ,When Tim Tebow found out he got cut by the Eagles he threw a fit...,0
post,3k6ady,2qh72,jokes,false,1441762692,https://old.reddit.com/r/Jokes/comments/3k6ady/a_boy_asks_his_jewish_father_for_50_dollars/,self.jokes,,"The father looked at his son and asked, ""40 dollars? What do you need 30 dollars for?""",A boy asks his Jewish father for 50 dollars...,9
post,3k692a,2qh72,jokes,false,1441762205,https://old.reddit.com/r/Jokes/comments/3k692a/pissing_in_the_snow/,self.jokes,,[deleted],Pissing in the snow...,3
post,3k68om,2qh72,jokes,false,1441762037,https://old.reddit.com/r/Jokes/comments/3k68om/what_do_you_call_nic_cage_when_hes_broke/,self.jokes,,"Nicolas (Nickle-less) Cage

stupidest thing I've ever come up with",What do you call Nic Cage when he's broke?,13
post,3k680b,2qh72,jokes,false,1441761776,https://old.reddit.com/r/Jokes/comments/3k680b/to_write_with_a_broken_pencil/,self.jokes,,[removed],to write with a broken pencil...,1
post,3k67lt,2qh72,jokes,false,1441761611,https://old.reddit.com/r/Jokes/comments/3k67lt/how_are_a_bad_mood_and_foreskin_alike/,self.jokes,,[deleted],How are a bad mood and foreskin alike?,0
post,3k675t,2qh72,jokes,false,1441761427,https://old.reddit.com/r/Jokes/comments/3k675t/go_fuck_yourself/,self.jokes,,"A kid walks up to his Grandpa and asks for a sip of his beer the Grandpa asks ""does you penis touch your asshole ?"" The kid says ""no"" The next day the kid asks for a sip of his Grandpa's beer and the Grandpa asks "" does your penis touch your asshole ? "" The kid says ""no"" So the next day the kid is eating a cookie and the Grandpa asks for a bite and the kid asks ""does your penis touch your butt ?"" the Grandpa says ""yes"" so the kid says ""go fuck yourself"".",Go fuck yourself,1
post,3k66an,2qh72,jokes,false,1441761085,https://old.reddit.com/r/Jokes/comments/3k66an/people_would_see_your_panties/,self.jokes,,"It was the first time for Jerry and his wife Agnes out of their little village, they headed to the city to attend the big festival.

When they reached there, the first thing that caught Agnes' eyes was the ferris wheel, she looked at her husband and asked him what it was, as she wanted to ride it, Jerry said ""it's called a ferris wheel, but you can't ride it, you're wearing a skirt and people would see your panties"" 

She kept nagging him for the next hour after each different ride saying she wants to try the ferris wheel and he kept replying ""People would see your panties"".

After another hour Jerry felt the need to go to the toilet, so he told his wife Agnes he's going to the toilet and he'd be back in 10 minutes, when he came back he looked for Agnes but couldn't find her, suddenly, she comes back running with a big smile on her face, he asks ""Where have you been?"" 

Agnes replies ""I rode the ferris wheel!""

Jerry says ""but people would see your panties!"" 

Agnes replies ""Don't worry, I took them off!""",People would see your panties!,5
post,3k666g,2qh72,jokes,false,1441761019,https://old.reddit.com/r/Jokes/comments/3k666g/a_couples_marriage_is_not_doing_so_well/,self.jokes,,[deleted],A couple's marriage is not doing so well...,1
post,3k6630,2qh72,jokes,false,1441760978,https://old.reddit.com/r/Jokes/comments/3k6630/whats_the_difference_between_broccoli_and_boogers/,self.jokes,,My son won't eat broccoli.,What's the difference between broccoli and boogers?,4
post,3k65zt,2qh72,jokes,false,1441760937,https://old.reddit.com/r/Jokes/comments/3k65zt/what_material_does_cayde6_use_to_repair_his_armor/,self.jokes,,"Nathan Filaments

( ͡° ͜ʖ ͡°)

X-Post from /r/DestinyTheGame",What material does Cayde-6 use to repair his armor after falling feet first into hell?,0
post,3k65ov,2qh72,jokes,false,1441760814,https://old.reddit.com/r/Jokes/comments/3k65ov/whats_a_racist_photographers_favorite_hobby/,self.jokes,,Crushing the blacks.,What's a racist photographer's favorite hobby?,0
post,3k6529,2qh72,jokes,false,1441760562,https://old.reddit.com/r/Jokes/comments/3k6529/one_day_superman_was_really_bored/,self.jokes,,"So he was flying around killing time. Suddenly he sees Wonder Woman spreadeagled naked on top of a tall building.

He has always fancied Wonder Woman so he thinks now's my chance as he swoops down and faster than a speeding bullet, does the business and then he flies off again.

A moment later Wonder Woman says ""what on earth was that?""

Then the Invisible Man climbs off her and says ""I don't know but my ass hurts a lot!""
",One day Superman was really bored...,10
post,3k63fr,2qh72,jokes,false,1441759961,https://old.reddit.com/r/Jokes/comments/3k63fr/three_nuns_die_and_end_up_at_the_gates_of_heaven/,self.jokes,,"Three nuns die and end up at the gates of Heaven.

St Peter says that before they can enter, they must first each answer a question.

To the first he asks ""who were the first humans?"" She says ""Adam and Eve"" and he lets her in.

To the second he asks ""where did they live?"" She says ""In the garden of Eden"" and she too is admitted.

Then he asks the third, ""what was the first thing Eve said to Adam?""

She replies ""My goodness that's a hard one"" - and he opens the gate and lets her in.",Three nuns die and end up at the gates of Heaven,0
post,3k6380,2qh72,jokes,false,1441759877,https://old.reddit.com/r/Jokes/comments/3k6380/mexican_word_of_the_day_nascar/,self.jokes,,Hey man that's a nascar..  Where'd you get it?,Mexican word of the day: nascar,0
post,3k632d,2qh72,jokes,false,1441759818,https://old.reddit.com/r/Jokes/comments/3k632d/the_bakery/,self.jokes,,"A guy named Rajesh works at a bakery in  Karachi, Pakistan. As a gopher, he is obligated to serve the baker. One day the baker says
""Raj, go and get me a bag of flour.""
Raj goes to get the bag and puts it on his head. Unfortunately the bag breaks and covers him from head to toe. Dejected, he walks back to the kitchen. 
""Oh my goodness Raj! What happened?""

""Well, I was carrying the bag of flour above my head and it broke so now I am going to go home and come back in 20 minutes.""

He walks out to the lobby where he meets the receptionist.
""Oh my goodness Raj! What happened?""

""Well, I was carrying the bag of flour above my head and it broke so now I am going to go home and come back in 20 minutes.""

Hopping on the same bus he rides everyday, the bus driver inquires:
""Oh my goodness Raj! What happened?""

""Well, I was carrying the bag of flour above my head and it broke so now I am going to go home and come back in 20 minutes.""

This happens a few more times on the way home. At the door to his home, he climbs the stairs, puts the key in the lock, and begins to twist when he is spotted by his neighbour.

""Oh my goodness, Raj! What happened?""

""GODDAMMIT! I have only been white for 10 minutes and already you fucking Pakis are getting on my nerves!""

Edit: changed the spelling of the racial slur so as to (oddly enough) be less offensive? Not sure how that works yet.",The Bakery,4
post,3k61py,2qh72,jokes,false,1441759311,https://old.reddit.com/r/Jokes/comments/3k61py/what_did_god_say_to_jesus/,self.jokes,,This lawn ain't gonna mow itself.,What did God say to Jesus?,0
post,3k60rh,2qh72,jokes,false,1441758934,https://old.reddit.com/r/Jokes/comments/3k60rh/how_do_you_turn_a_gay_man_straight/,self.jokes,,Give him a beard,How do you turn a gay man straight?,0
post,3k60q6,2qh72,jokes,false,1441758919,https://old.reddit.com/r/Jokes/comments/3k60q6/i_went_to_my_marriage_counsellor_today_nsfw/,self.jokes,,"I told him I wasn't sexually attracted to my wife anymore, He asked why I said she's just too lose, and I can't feel anything I just don't enjoy it as much as i used too. He suggested to me why don't i try the other hole? So i replied no way! she can get pregnant from that one.
",I went to my marriage counsellor today [NSFW],1
post,3k6067,2qh72,jokes,false,1441758664,https://old.reddit.com/r/Jokes/comments/3k6067/how_do_white_supremacists_celebrate_their/,self.jokes,,[deleted],How do white supremacists celebrate their birthdays?,1
post,3k5zw1,2qh72,jokes,false,1441758535,https://old.reddit.com/r/Jokes/comments/3k5zw1/how_many_licks_does_it_take_to_pop_a_cherry/,self.jokes,,[deleted],How many licks does it take to pop a cherry?,0
post,3k5zjc,2qh72,jokes,false,1441758394,https://old.reddit.com/r/Jokes/comments/3k5zjc/what_do_you_call_a_midget_mexican/,self.jokes,,A little Juan.,What do you call a midget Mexican?,13
post,3k5z1t,2qh72,jokes,false,1441758218,https://old.reddit.com/r/Jokes/comments/3k5z1t/shetoldme/,self.jokes,,[removed],#SheToldMe 01001000011000010111001101101000011101000110000101100111,1
post,3k5yno,2qh72,jokes,false,1441758073,https://old.reddit.com/r/Jokes/comments/3k5yno/who_would_guess_that_people_will_fight_to_get/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k5yno/who_would_guess_that_people_will_fight_to_get/,,Who would guess that people will fight to get into trains heading for German camps.,3
post,3k5xy4,2qh72,jokes,false,1441757813,https://old.reddit.com/r/Jokes/comments/3k5xy4/the_man_with_the_25_inch_penis/,self.jokes,,"A man who had a 25 inch long penis went to his doctor to complain that he was having a problem with this rather massive instrument and has had more than one complaint. ""Doctor,"" he asked, in total frustration, ""is there anything you can do for me?"" The doctor replies, ""Medically son, there is nothing I can do. But, I do know this witch who may be able to help you."" So the doctor gives him directions to the witch.

The man calls upon the witch and relays his story. ""Witch, my penis is 25 inches long and I need help. Can anything be done to help me? You are my last hope!"" The witch stares in amazement, scratches her head, and then replies, ""I think I may be able to help you. Do this. Go deep into the forest. You will find a pond. In this pond, you will find a frog sitting on a log. This frog has magic. You say to frog, will you marry me? When the frog says no, you will find five inches less to your problem."" The man's face lit up and he dashed off into the forest. He called out to the frog, ""Will you marry me?""

The frog looked at him dejectedly and replied, ""NO."" The man looked down and suddenly his penis was 5 inches shorter. ""WOW,"" he screamed out loud, ""This is great!!"" But at 20 inches it was still too long, so he asked the frog again. ""Frog, will you marry me?"" the guy shouted. The frog rolled its eyes back in its head and screamed back, ""NO!"" The man felt another twitch in his penis, looked down, and it was another 5 inches shorter. The man laughed, ""This is fantastic."" He looked down at his penis again, 15 inches long, and reflected for a moment Fifteen inches is still a monster, just a little less would be ideal.

Grinning, he looked across the pond and yelled out, ""Frog will you marry me?"" The frog looked back across pond shaking its head, ""How many times do I have to tell you? NO, NO, NO!!""
",The man with the 25 inch penis,12
post,3k5x0x,2qh72,jokes,false,1441757466,https://old.reddit.com/r/Jokes/comments/3k5x0x/why_do_you_call_how_do_you/,self.jokes,,[removed],Why do you call? How do you? 0101100101101111001000000100110101101111011011010110110101100001,1
post,3k5x0g,2qh72,jokes,false,1441757463,https://old.reddit.com/r/Jokes/comments/3k5x0g/how_to_prove_jokeexplainbot_is_actually_a_human/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k5x0g/how_to_prove_jokeexplainbot_is_actually_a_human/,,How to prove JokeExplainBot is actually a human?,1
post,3k5wt4,2qh72,jokes,false,1441757378,https://old.reddit.com/r/Jokes/comments/3k5wt4/jewish_joke_about_warm_weather/,self.jokes,,"אחי היה לי כלכך חם שהבטחתי שאם יציעו לי להתנצר בזה הרגע אני אעשה את זה רק בשביל ההטבלה.

Dude. It was so hot, I swear that I'd convert to Christianity for the Baptism.",Jewish Joke About Warm Weather,5
post,3k5wsy,2qh72,jokes,false,1441757376,https://old.reddit.com/r/Jokes/comments/3k5wsy/why_does_a_man_refuse_to_listen_to_his_front_seat/,self.jokes,,[deleted],Why does a man refuse to listen to his front seat passenger when he is lost?,5
post,3k5wlr,2qh72,jokes,false,1441757302,https://old.reddit.com/r/Jokes/comments/3k5wlr/what_did_the_pink_panther_say_when_he_stepped_on/,self.jokes,,"Dead ant 
Dead ant 
Dead ant dead ant dead ant
Dead ant dead annnnnnt 
Dead ant",What did the Pink Panther say when he stepped on an ant?,4
post,3k5u0c,2qh72,jokes,false,1441756304,https://old.reddit.com/r/Jokes/comments/3k5u0c/you_have_a_dime_in_one_hand_and_a_nickel_in_the/,self.jokes,,Broke.,You have a dime in one hand and a nickel in the other. What are you?,7
post,3k5tki,2qh72,jokes,false,1441756121,https://old.reddit.com/r/Jokes/comments/3k5tki/how_many_dead_whores_does_it_take_to_change_a/,self.jokes,,"More than three, I still can't reach it.",How many dead whores does it take to change a light bulb?,48
post,3k5thm,2qh72,jokes,false,1441756088,https://old.reddit.com/r/Jokes/comments/3k5thm/whats_the_difference_between_bigfoot_and_a/,self.jokes,,Bigfoot is occasionally sighted,What's the difference between Bigfoot and a Mexican with a beard?,0
post,3k5t74,2qh72,jokes,false,1441755982,https://old.reddit.com/r/Jokes/comments/3k5t74/there_are_three_kinds_of_people/,self.jokes,,"The ones that can count, and the ones that can't.",There are three kinds of people,2
post,3k5s87,2qh72,jokes,false,1441755597,https://old.reddit.com/r/Jokes/comments/3k5s87/whats_the_best_way_to_kill_a_bug/,self.jokes,,Just bug him to death.,What's the best way to kill a bug?,3
post,3k5rzg,2qh72,jokes,false,1441755510,https://old.reddit.com/r/Jokes/comments/3k5rzg/whats_the_difference_between_here_and_there/,self.jokes,,"When you're right the whole room shouts ""Here, here!"" But when you're wrong one person pats you on the back and says ""There, there.""",What's the difference between Here and There?,6
post,3k5rdd,2qh72,jokes,false,1441755261,https://old.reddit.com/r/Jokes/comments/3k5rdd/i_would_start_an_auto_cannibalistic_society/,self.jokes,,[deleted],I would start an auto cannibalistic society...,1
post,3k5qk6,2qh72,jokes,false,1441754928,https://old.reddit.com/r/Jokes/comments/3k5qk6/what_did_the_dog_say_to_the_fireman/,self.jokes,,The roof is on fire.,What did the dog say to the fireman?,0
post,3k5q9j,2qh72,jokes,false,1441754807,https://old.reddit.com/r/Jokes/comments/3k5q9j/there_are_six_american_flags_on_the_moon/,self.jokes,,"Five of them are still standing. Due to the strong UV radiation, they are all completely white by now.

So it looks like the French landed there.",There are six American flags on the Moon.,84
post,3k5oqk,2qh72,jokes,false,1441754203,https://old.reddit.com/r/Jokes/comments/3k5oqk/my_son_dropped_this_gem_on_me/,self.jokes,,"Son: Dad what's a cow plus 2 say?

Me: Cow cow?

Son: Twwoooooooooo",My son dropped this gem on me,1
post,3k5oq9,2qh72,jokes,false,1441754200,https://old.reddit.com/r/Jokes/comments/3k5oq9/a_mexican_walked_into_a_polish_store_and_greeted/,self.jokes,,"He was handed a sausage.

Edit: Ok I will walk myself out...",A Mexican walked into a Polish store and greeted every one.,0
post,3k5omn,2qh72,jokes,false,1441754169,https://old.reddit.com/r/Jokes/comments/3k5omn/dating_in_your_30s_is_like_looking_for_a_parking/,self.jokes,,The good ones are all taken.  The rest are either handicapped or too far away.,Dating in your 30s is like looking for a parking spot...,7113
post,3k5o9d,2qh72,jokes,false,1441754042,https://old.reddit.com/r/Jokes/comments/3k5o9d/two_balloons_are_floating_through_the_desert/,self.jokes,,[deleted],Two balloons are floating through the desert...,0
post,3k5nas,2qh72,jokes,false,1441753637,https://old.reddit.com/r/Jokes/comments/3k5nas/a_jew_a_catholic_and_a_mormon_are_drinking/,self.jokes,,"The Jew boasts about his fertility

""I have 4 sons; one more and I'll have a basketball team!""

""That's nothing,"" says the Catholic, ""I have 10 sons! I almost have a football team!""

The Jew and Catholic looked expectantly at the Mormon. ""Well?""

""I have 17 wives. I almost have a golf course!""","A Jew, a Catholic, and a Mormon are drinking together.",648
post,3k5n14,2qh72,jokes,false,1441753558,https://old.reddit.com/r/Jokes/comments/3k5n14/q_do_you_think_id_be_a_good_parent/,self.jokes,,[deleted],"Q: ""Do you think I'd be a good parent?""",1
post,3k5mmi,2qh72,jokes,false,1441753400,https://old.reddit.com/r/Jokes/comments/3k5mmi/friends_wife_told_me_a_joke/,self.jokes,,[deleted],Friends wife told me a joke,0
post,3k5lfq,2qh72,jokes,false,1441752961,https://old.reddit.com/r/Jokes/comments/3k5lfq/an_elderly_couple_file_for_divorce/,self.jokes,,"... After 60 years of marriage. The lawyer they meet with prepares all the paperwork but stops before handing it to the couple to sign and asks;

""By all means I can let you do this, but please let me know why? Why after over half a century of happy marriage would you want to end it now? What could ruin such a long streak of love?""

""Well,"" replies the wife, ""we wanted to wait until the kids were dead."" ",An elderly couple file for divorce...,3
post,3k5ky2,2qh72,jokes,false,1441752762,https://old.reddit.com/r/Jokes/comments/3k5ky2/an_elementary_teacher_told_her_students_that_if/,self.jokes,,"The teacher asked, ""Who said 'A house divided against itself cannot stand'?"" 
Susan in the front raised her hand and said ""Abraham Lincoln"" and she was allowed to leave.
The teacher then asked, ""Who said 'Ask not what your country can do for you, but what you can do for your country'?""
Abby, who was also sitting in the front, raised her hand and said ""John F Kennedy"" and she was allowed to leave.
This whole time John, who was sitting in the back and really wanted to go home, had known all the right answers but was not getting called on because he was sitting in the back. He muttered to himself, ""If only those girls had kept quiet, I wouldn't have to be in this situation."" 
""Who said that?"" The teacher called out.
""Bill Clinton!"" Shouted John. He gathered his stuff and went home.",An elementary teacher told her students that if they could answer the questions correctly they would be dismissed from class.,2
post,3k5k0b,2qh72,jokes,false,1441752413,https://old.reddit.com/r/Jokes/comments/3k5k0b/have_you_heard_of_the_new_pencils_theyre/,self.jokes,,[deleted],Have you heard of the new pencils they're developing with no lead?,0
post,3k5it2,2qh72,jokes,false,1441751965,https://old.reddit.com/r/Jokes/comments/3k5it2/sodium_sodium_sodium_sodium_sodium_sodium_sodium/,self.jokes,,[deleted],Sodium Sodium Sodium Sodium Sodium Sodium Sodium Sodium Sodium Boron Argon Titanium Manganese!,0
post,3k5isb,2qh72,jokes,false,1441751958,https://old.reddit.com/r/Jokes/comments/3k5isb/adam_sandler/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k5isb/adam_sandler/,,Adam Sandler,0
post,3k5icd,2qh72,jokes,false,1441751799,https://old.reddit.com/r/Jokes/comments/3k5icd/how_do_you_think_the_unthinkable/,self.jokes,,With an Itheberg,How do you think the unthinkable?,80
post,3k5gvx,2qh72,jokes,false,1441751276,https://old.reddit.com/r/Jokes/comments/3k5gvx/a_man_was_caught_peeing_in_public_by_a_police/,self.jokes,,"""Urine trouble now.""",A man was caught peeing in public by a police officer. The cop's only reaction was...,5
post,3k5fts,2qh72,jokes,false,1441750882,https://old.reddit.com/r/Jokes/comments/3k5fts/my_mexican_friend_told_me_he_is_far_sided_i_said/,self.jokes,,"to which he replied

&gt;""No, I *quinceanera*""","My mexican friend told me he is far sided, I said so does that mean you cant see far away?",0
post,3k5frv,2qh72,jokes,false,1441750859,https://old.reddit.com/r/Jokes/comments/3k5frv/john_mcafees_doing_paper_work_to_become_president/,self.jokes,,Time for America to become bloated and slow...,John McAfee's doing paper work to become president...,0
post,3k5esu,2qh72,jokes,false,1441750503,https://old.reddit.com/r/Jokes/comments/3k5esu/how_can_you_tell_a_mechanic_just_had_sex/,self.jokes,,Two of his fingers are clean.,How can you tell a mechanic just had sex?,598
post,3k5dd6,2qh72,jokes,false,1441749907,https://old.reddit.com/r/Jokes/comments/3k5dd6/fishing/,self.jokes,,"A local sheriff received an anonymous tip that there was a young man fishing at the pond without a license. He decides to check it out, and, arriving at the pond, he spots two teenagers fishing at the shore. As he is approaching the pair, one of them looks up, sees the sheriff, and takes off at a sprint. He gives chase, trailing him for about a quarter-mile, at which point the young man is out of breath. 
     The sheriff grabs him and says, panting, ""Let me see your fishing license."" The teenager pulls out his license and hands it to him. ""Why'd you run away from me if you have a license? You weren't doing anything wrong,"" the policeman gasps, still exhausted.
      Suddenly, a grin appears on the young man's face. ""I have my license,"" he explained, ""but my buddy back there doesnt!""",Fishing,14
post,3k5d2t,2qh72,jokes,false,1441749790,https://old.reddit.com/r/Jokes/comments/3k5d2t/what_do_you_call_a_bird_with_a_teacup_on_its_head/,self.jokes,,[deleted],What do you call a bird with a teacup on its head?,1
post,3k5cpn,2qh72,jokes,false,1441749642,https://old.reddit.com/r/Jokes/comments/3k5cpn/what_did_the_conceited_man_say_while_he_stood_on/,self.jokes,,The earth revolves around me.,What did the conceited man say while he stood on the north pole?,0
post,3k5btp,2qh72,jokes,false,1441749304,https://old.reddit.com/r/Jokes/comments/3k5btp/they_told_me_i_had_type_a_blood/,self.jokes,,But it was a type O.,They told me i had type A blood.,313
post,3k5b9a,2qh72,jokes,false,1441748992,https://old.reddit.com/r/Jokes/comments/3k5b9a/how_to_know_shes_the_one/,self.jokes,,"Jerk off twice and if you still wanna jerk off, then She is.",How to know she's the one?,0
post,3k5avq,2qh72,jokes,false,1441748815,https://old.reddit.com/r/Jokes/comments/3k5avq/i_heard_the_problems_in_syria_are_because_of_some/,self.jokes,,[deleted],I heard the problems in Syria are because of some...,0
post,3k59y6,2qh72,jokes,false,1441748400,https://old.reddit.com/r/Jokes/comments/3k59y6/can_i_have_some_of_that_well/,self.jokes,,"An old man takes his grandson to the bar. The grandfather orders a whiskey, takes a swig, then puts it down.

The kid asks, ""Hey grandpa, can I have some of that?""

Grandpa replies, ""Does the tip of your dick reach the cheeks of your ass?""

""Nope.""

""Well there's your answer.""

After a little while of drinking, the grandfather pulls out a pack of cigarettes and lights one up.

The kids asks, ""Hey grandpa, can I get one of those?""

""Does the tip of your dick reach the cheeks of your ass?""

""Nope.""

""Well there's your answer.""

So after a little while they get tired and pack up to go home. On the way home they stop at a little store, and each buys a lottery ticket. Grandpa scratches his and wins nothing.

The grandson scratches his and wins $5,000.

Grandpa asks, ""Hey kid, can I have some of that?""

""Does the tip of your dick reach the cheeks of your ass?""

""Sure does.""

""Well then you can go fuck yourself cuz you ain't gettin' none of this.""",Can I have some of that? Well...,5
post,3k595u,2qh72,jokes,false,1441748076,https://old.reddit.com/r/Jokes/comments/3k595u/how_often_do_i_make_jokes_about_chemistry/,self.jokes,,Periodically.,How often do i make jokes about chemistry?,38
post,3k57pv,2qh72,jokes,false,1441747490,https://old.reddit.com/r/Jokes/comments/3k57pv/can_i_get_have_of_that_well/,self.jokes,,[deleted],Can I get have of that? Well...,1
post,3k56lz,2qh72,jokes,false,1441747011,https://old.reddit.com/r/Jokes/comments/3k56lz/joke_from_my_niece/,self.jokes,,"Her: Why did the chicken cross the road?
 Me: Why?
 Her: To get to the ugly guy's house. 
Me:??? 
Her: Knock knock
 Me: Who's there? 
Her: It's the chicken!",Joke From My Niece,10
post,3k560l,2qh72,jokes,false,1441746753,https://old.reddit.com/r/Jokes/comments/3k560l/how_to_piss_off_the_jokeexplainbot/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k560l/how_to_piss_off_the_jokeexplainbot/,,How to piss off the JokeExplainBot?,1
post,3k55ui,2qh72,jokes,false,1441746674,https://old.reddit.com/r/Jokes/comments/3k55ui/a_roman_man_walks_into_a_bar_and_holds_up_two/,self.jokes,,[deleted],A roman man walks into a bar and holds up two fingers,5
post,3k55a9,2qh72,jokes,false,1441746427,https://old.reddit.com/r/Jokes/comments/3k55a9/what_do_you_call_it_when_stevie_wonder_and_ray/,self.jokes,,Endless Love,What do you call it when Stevie Wonder and Ray Charles play tennis?,121
post,3k555i,2qh72,jokes,false,1441746376,https://old.reddit.com/r/Jokes/comments/3k555i/the_joneses_and_the_whitneys_decide_to_go_swinging/,self.jokes,,"They go to a cabin motel, each couple gets a cabin, and after a good supper in a nearby restaurant and a camp fire, they all go to bed in their cabins.

The next morning, Mr Jones wakes up and says: ""Hmmm, that was a good night. Let's go see how the wives are doing""...",The Joneses and the Whitneys decide to go swinging...,0
post,3k554i,2qh72,jokes,false,1441746365,https://old.reddit.com/r/Jokes/comments/3k554i/kim_daviss_daughter_was_fired_by_the_spca/,self.jokes,,She wouldn't feed the strays,Kim Davis's Daughter was Fired by the SPCA,5
post,3k54ls,2qh72,jokes,false,1441746153,https://old.reddit.com/r/Jokes/comments/3k54ls/question_about_god/,self.jokes,,if god can do anything can he do nothing?,question about god?,0
post,3k54ai,2qh72,jokes,false,1441746034,https://old.reddit.com/r/Jokes/comments/3k54ai/a_young_boy_was_riding_with_his_new_bike_and_goes/,self.jokes,,[deleted],A young boy was riding with his new bike and goes to talk with a mounted policeman.,0
post,3k53et,2qh72,jokes,false,1441745667,https://old.reddit.com/r/Jokes/comments/3k53et/a_friend_of_mine_died_in_the_middle_of_an_orgy/,self.jokes,,I'm glad he spent his final moments surrounded by his family. ,A friend of mine died in the middle of an orgy,3
post,3k52j2,2qh72,jokes,false,1441745287,https://old.reddit.com/r/Jokes/comments/3k52j2/knock_knock_whos_there_911/,self.jokes,,"Knock knock?
Who’s there?
9/11.
9/11 who?
You said you would never forget… :(
",Knock knock? Who’s there? 9/11,64
post,3k528x,2qh72,jokes,false,1441745173,https://old.reddit.com/r/Jokes/comments/3k528x/what_do_you_call_a_terrorists_girlfriend/,self.jokes,,"A Guantanamo Bae


Thought of this one earlier and just had to share",What do you call a terrorist's girlfriend?,1749
post,3k50hf,2qh72,jokes,false,1441744391,https://old.reddit.com/r/Jokes/comments/3k50hf/johnny_asked_to_sam/,self.jokes,,"Johnny asked to Sam what they will do that night.
Sam said “we will flip a coin
Then Johnny said “If it comes head, we will go for movies. If tails, we will play cards, if it stands on edge, we will study",Johnny asked to Sam,0
post,3k5092,2qh72,jokes,false,1441744304,https://old.reddit.com/r/Jokes/comments/3k5092/a_young_couple_goes_to_a_party/,self.jokes,,"The young lady, being a bit of a princess, tells the young man that he must first sample all of the drinks, bring her the best one and then tell her a joke to start the party. The young man samples all of the drinks and returns with a tequila sunrise. 
""What about my joke?""
""Ok,"" he replies, ""a man walks in to a bar, has a drink and goes home.""
""That's the joke?""
""There is no punch line!!!"" She exclaims.
""And there won't be, the punch here tastes like shit.""",A young couple goes to a party.,2
post,3k4zyr,2qh72,jokes,false,1441744208,https://old.reddit.com/r/Jokes/comments/3k4zyr/just_remember_youre_unique/,self.jokes,,Just like everyone else.,"Just remember, you're unique.",0
post,3k4zn6,2qh72,jokes,false,1441744017,https://old.reddit.com/r/Jokes/comments/3k4zn6/whats_the_difference_between_firewood_and_a_jew/,self.jokes,,The firewood ain't been turned into ash yet.,What's the difference between firewood and a jew?,0
post,3k4yy2,2qh72,jokes,false,1441743708,https://old.reddit.com/r/Jokes/comments/3k4yy2/nsfw_we_all_want_something/,self.jokes,,"White people: legalize gay marriage!!
Black people: legalize weed!!
Mexicans: legalize us!!",(NSFW) we all want something...,0
post,3k4yw1,2qh72,jokes,false,1441743686,https://old.reddit.com/r/Jokes/comments/3k4yw1/my_wife_got_mad_at_me_for_starting_another/,self.jokes,,"I said, ""don't worry, it'll be over soon.""",My wife got mad at me for starting another British TV series...,4
post,3k4ykl,2qh72,jokes,false,1441743561,https://old.reddit.com/r/Jokes/comments/3k4ykl/if_bernie_sanders_gets_elected_they_should_rename/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k4ykl/if_bernie_sanders_gets_elected_they_should_rename/,,"If Bernie Sanders gets elected, they should rename the White House the ""Sand Castle"".",0
post,3k4yhk,2qh72,jokes,false,1441743529,https://old.reddit.com/r/Jokes/comments/3k4yhk/two_guys_were_picked_up_by_the_cops/,self.jokes,,[deleted],Two guys were picked up by the cops!,2
post,3k4xse,2qh72,jokes,false,1441743249,https://old.reddit.com/r/Jokes/comments/3k4xse/on_a_traffic_light_green_means_go_yellow_means/,self.jokes,,"But on a banana it's just the opposite. Green means hold on, yellow means go ahead, and red means where the fuck did you get that banana at?","On a traffic light green means go, yellow means yield and red means stop.",3
post,3k4w2y,2qh72,jokes,false,1441742543,https://old.reddit.com/r/Jokes/comments/3k4w2y/a_boss_said_to_his_secretary_i_want_to_have_sex/,self.jokes,,"She thought for a moment then called her boyfriend and told him the story.  Her boyfriend then said to her, do it but ""Ask him for $2000, pick up the money very fast he wouldn't even have enough time to undressed himself.""  So she agrees. Half an hour goes by, the boyfriend decides to call girlfriend, he asks, what happened?  She responds, ""The Bastard used coins I'm still picking and he is still fucking!","A boss said to his secretary I want to have SEX with you I will make it very fast. I'll throw $1000 on the floor, by the time you bend down to pick it I'll be done.",11
post,3k4tnt,2qh72,jokes,false,1441741597,https://old.reddit.com/r/Jokes/comments/3k4tnt/its_so_rude_when_someones_phone_goes_off_in_class/,self.jokes,,Some of us are trying to sleep.,It's so rude when someone's phone goes off in class.,489
post,3k4sej,2qh72,jokes,false,1441741054,https://old.reddit.com/r/Jokes/comments/3k4sej/knock_knock/,self.jokes,,"""Who's there?""

""Allah!""

""Allah who?""

""ALLAHU AKBAR!!""","""Knock Knock!""",0
post,3k4s0p,2qh72,jokes,false,1441740892,https://old.reddit.com/r/Jokes/comments/3k4s0p/husband_wife/,self.jokes,,[deleted],husband wife,0
post,3k4r2u,2qh72,jokes,false,1441740511,https://old.reddit.com/r/Jokes/comments/3k4r2u/i_received_an_email_from_google/,self.jokes,,"It said, ""At Google Earth we can read maps backwards "" I thought, ""That's just spam."" ",I received an email from Google,1618
post,3k4o64,2qh72,jokes,false,1441739304,https://old.reddit.com/r/Jokes/comments/3k4o64/wes_craven_died/,self.jokes,,"Well that sucks, I sure wes craven another scary movie...",Wes Craven died?,0
post,3k4o41,2qh72,jokes,false,1441739278,https://old.reddit.com/r/Jokes/comments/3k4o41/did_you_guys_hear_about_the_homeopath_who_forgot/,self.jokes,,He died of an overdose.,Did you guys hear about the homeopath who forgot to take his meds?,2
post,3k4nwl,2qh72,jokes,false,1441739200,https://old.reddit.com/r/Jokes/comments/3k4nwl/dyslexic_man/,self.jokes,,[deleted],Dyslexic man,3
post,3k4nl6,2qh72,jokes,false,1441739074,https://old.reddit.com/r/Jokes/comments/3k4nl6/my_teacher_told_me_that_my_test_results_were/,self.jokes,,"Me: Really? They're that good? 

Teacher: No they're utterly terrible but we can absolutely get them re-marked by the exam board and turn that F- into an F. ","My teacher told me that my test results were ""absolutely remarkable""...",0
post,3k4mde,2qh72,jokes,false,1441738576,https://old.reddit.com/r/Jokes/comments/3k4mde/she_takes_up_two_jokes/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k4mde/she_takes_up_two_jokes/,,She takes up two jokes,0
post,3k4lop,2qh72,jokes,false,1441738321,https://old.reddit.com/r/Jokes/comments/3k4lop/whats_long_brown_and_sticky/,self.jokes,,A stick,"What's long, brown, and sticky?",0
post,3k4ln1,2qh72,jokes,false,1441738302,https://old.reddit.com/r/Jokes/comments/3k4ln1/what_is_the_best_cabinet_post_for_donald_trump/,self.jokes,,"Secretary of 'De-Fence""",What is the best Cabinet post for Donald Trump?,0
post,3k4lll,2qh72,jokes,false,1441738284,https://old.reddit.com/r/Jokes/comments/3k4lll/what_genre_of_porn_does_the_pope_watch/,self.jokes,,[deleted],What genre of porn does the Pope watch?,1
post,3k4l59,2qh72,jokes,false,1441738109,https://old.reddit.com/r/Jokes/comments/3k4l59/what_is_it_called_when_more_than_one_hundred/,self.jokes,,[deleted],What is it called when more than one hundred people agree with you on Reddit?,0
post,3k4kib,2qh72,jokes,false,1441737853,https://old.reddit.com/r/Jokes/comments/3k4kib/i_went_for_a_meal_at_my_local_chinese_restaurant/,self.jokes,,...I don't even like Chinese food but I thought I'd check it out because people keep telling me that God works there. ,"I went for a meal at my local Chinese restaurant ""Mysterious Ways"" yesterday...",0
post,3k4ki5,2qh72,jokes,false,1441737852,https://old.reddit.com/r/Jokes/comments/3k4ki5/yo_momma_so_fat/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k4ki5/yo_momma_so_fat/,,Yo momma so fat,0
post,3k4kfd,2qh72,jokes,false,1441737819,https://old.reddit.com/r/Jokes/comments/3k4kfd/what_do_you_call_a_tightfisted_wookie/,self.jokes,,Jewbacca,What do you call a tight-fisted Wookie?,0
post,3k4jjd,2qh72,jokes,false,1441737462,https://old.reddit.com/r/Jokes/comments/3k4jjd/whats_soulja_boys_favorite_letter_in_the_cyrillic/,self.jokes,,[deleted],What's Soulja Boy's favorite letter in the Cyrillic alphabet?,0
post,3k4ims,2qh72,jokes,false,1441737093,https://old.reddit.com/r/Jokes/comments/3k4ims/you_dont_need_a_parachute_to_go_skydiving/,self.jokes,,..You need a parachute to go skydiving twice.,You don’t need a parachute to go skydiving..,11
post,3k4i7g,2qh72,jokes,false,1441736914,https://old.reddit.com/r/Jokes/comments/3k4i7g/that_stupid_guy/,self.jokes,,I have stupid friends gotta admit.But i have a stupid one. Yesterday he asked me did anybody die and survive??!?!?!??,That stupid guy,0
post,3k4hfo,2qh72,jokes,false,1441736588,https://old.reddit.com/r/Jokes/comments/3k4hfo/tifu_misinterpreting_an_acronym/,self.jokes,,[deleted],TIFU misinterpreting an acronym.,0
post,3k4h3f,2qh72,jokes,false,1441736466,https://old.reddit.com/r/Jokes/comments/3k4h3f/why_did_the_chicken_fall_in_the_well/,self.jokes,,Because he couldn't see that well!,Why did the chicken fall in the well?,24
post,3k4gih,2qh72,jokes,false,1441736215,https://old.reddit.com/r/Jokes/comments/3k4gih/racist_jokes/,self.jokes,,Go!,Racist jokes...,0
post,3k4f0o,2qh72,jokes,false,1441735625,https://old.reddit.com/r/Jokes/comments/3k4f0o/damn_i_burnt_one/,self.jokes,,"What did God say when he made the first black man? 

""Damn, I burnt one."" ","Damn, I burnt one.",0
post,3k4eo3,2qh72,jokes,false,1441735490,https://old.reddit.com/r/Jokes/comments/3k4eo3/what_do_you_call_a_mexican_midget/,self.jokes,,A paragraph because he's not a full ese.,What do you call a Mexican midget?,1
post,3k4doe,2qh72,jokes,false,1441735091,https://old.reddit.com/r/Jokes/comments/3k4doe/a_chicken_walks_into_a_library/,self.jokes,,"...and goes up to the circulation desk. ""Bok!"" he says. The clerk thought for a moment and then said, ""Oh! You want a book!"" So he gives the chicken a book and the chicken walks out.

A few hours later the chicken comes back and says, ""Bok bok!"" The clerk thinks to himself that that was a little fast to read a book, but checks out two more for the chicken and the chicken walks out. 

A third time the chicken comes in and wails, ""Bok, bok, BOK!"" Thoroughly confused, the clerk checks out three new books for the chicken but decides to follow him instead. The chicken walks into the woods, over a hill, and down to a pond, with the clerk following at a distance. The chicken walks to the water's edge and drops the books in front of a frog. The frog looks at the first book at says, ""reddit.""",A chicken walks into a library...,152
post,3k4btm,2qh72,jokes,false,1441734356,https://old.reddit.com/r/Jokes/comments/3k4btm/mike_tyson_mysteries_is_on_netflix_now/,self.jokes,,Episode 1: case of the missing ear.,Mike Tyson Mysteries is on Netflix now...,0
post,3k4boq,2qh72,jokes,false,1441734306,https://old.reddit.com/r/Jokes/comments/3k4boq/what_happens_when_a_spanish_person_and_a_french/,self.jokes,,They give birth to an Andorran.,What happens when a Spanish person and a French person fuck?,0
post,3k4bdn,2qh72,jokes,false,1441734198,https://old.reddit.com/r/Jokes/comments/3k4bdn/have_a_coke_and_a_smile/,self.jokes,,"I opened up a can of Coke, and on the side it said: ""Share a Coke with your Soulmate."" So, I put the can in my right hand.",Have a Coke and a smile!,1
post,3k4b6z,2qh72,jokes,false,1441734121,https://old.reddit.com/r/Jokes/comments/3k4b6z/you_get_out_of_life_what_you_put_in_to_it/,self.jokes,,[removed],You get out of life what you put in to it,1
post,3k4a6e,2qh72,jokes,false,1441733706,https://old.reddit.com/r/Jokes/comments/3k4a6e/an_austrian_drunk_is_passing_by_a_cemetery/,self.jokes,,"An Austrian drunk is passing by a cemetery, when he hears music, following the music, he finds its coming from a grave, frightened, he begins to run away and bumps into a policeman. 

'Vere are you going at zis hour?' asks the policeman, 

'Entschuldigung, I've been celebrating, I was walking past ze cemetery, when I heard music' 

'Music? In ze cemetery?'

'Ja, but I'm drunk so might not be'

'Lets check it out.'

The cop hears the music too, and decides to go to the nearby church and fetch a priest. 

The priest arrives and listens ' Ah! Zat is Herr Mozart's 5th symphony... but it is being played backvords, and zere, it is now the 4th, also being played backvords....' 

The priest finally realizes ' Ah! Nothing to worry, it is just Herr Mozart decomposing' ",An austrian drunk is passing by a cemetery...,9
post,3k49z7,2qh72,jokes,false,1441733625,https://old.reddit.com/r/Jokes/comments/3k49z7/why_do_elephants_drink_so_much/,self.jokes,,To try to forget!,Why do elephants drink so much?,0
post,3k49qm,2qh72,jokes,false,1441733526,https://old.reddit.com/r/Jokes/comments/3k49qm/freudian_slip/,self.jokes,,[deleted],Freudian slip:,0
post,3k48iy,2qh72,jokes,false,1441733034,https://old.reddit.com/r/Jokes/comments/3k48iy/drunk_welsh_man_walks_into_a_bar/,self.jokes,,"A drunk welsh man walks into a bar. How many women are pregnant at the end of the night?   None, but I wouldn't eat the lamb!
",Drunk Welsh man walks into a bar,3
post,3k47y4,2qh72,jokes,false,1441732806,https://old.reddit.com/r/Jokes/comments/3k47y4/a_boat_in_the_atlantic_ocean_was_starting_to_sink/,self.jokes,,"... The captain gathered everyone and said ""OK everyone, it looks like we are going down, does anyone know how to pray?"" One of the ships crew members sitting in the back raises his hand and Hays ""yes captain I know how to pray."" The captain responds ""OK well you start praying and everyone else put a life jacket on, we're short one jacket.""

Another joke from my 95 year old grandpa. ",A boat in the Atlantic ocean was starting to sink...,47
post,3k47uj,2qh72,jokes,false,1441732767,https://old.reddit.com/r/Jokes/comments/3k47uj/my_cheap_boss/,self.jokes,,Talks so much shit. I guess its hard to defecate when you're major tight ass.,My cheap boss...,0
post,3k47dg,2qh72,jokes,false,1441732573,https://old.reddit.com/r/Jokes/comments/3k47dg/two_women_talking/,self.jokes,,"""Last night my man gave me a nice bouquet of flowers and took me to the fanciest restaurant to celebrate our anniversary. I thought to myself, girl, you'll have to spread those legs when we get back home!""

""Didn't you have at least a vase or something?""",Two women talking,1
post,3k473z,2qh72,jokes,false,1441732479,https://old.reddit.com/r/Jokes/comments/3k473z/this_is_the_punchline/,self.jokes,,[deleted],This is the punchline.,0
post,3k45w7,2qh72,jokes,false,1441732006,https://old.reddit.com/r/Jokes/comments/3k45w7/what_is_laziness_logical_answer/,self.jokes,,It is the Art of Taking Rest Before Getting Tired.,What is Laziness? Logical Answer,0
post,3k45w3,2qh72,jokes,false,1441732004,https://old.reddit.com/r/Jokes/comments/3k45w3/how_did_the_underage_mathematician_get_drunk/,self.jokes,,He put his root beer in a square glass,How did the underage mathematician get drunk?,220
post,3k44lr,2qh72,jokes,false,1441731536,https://old.reddit.com/r/Jokes/comments/3k44lr/how_many_jews_does_it_take_to_kill_jesus/,self.jokes,,You can't kill a myth.,How many Jews does it take to kill Jesus?,0
post,3k43ej,2qh72,jokes,false,1441731073,https://old.reddit.com/r/Jokes/comments/3k43ej/how_do_you_make_a_baby_cry_twice/,self.jokes,,You rub your bloody dick on their teddy bear. ,How do you make a baby cry twice?,0
post,3k41qm,2qh72,jokes,false,1441730405,https://old.reddit.com/r/Jokes/comments/3k41qm/a_little_boy_in_a_very_catholic_school_sharted/,self.jokes,,"The teacher promptly hands him a note and says that he has been fined 75 pence for unwarranted behaviour. She further explains that the little boy has to pay 50 cents for sharting and a quarter for peeing his pants.  
The little boy took the note, read it, but seemed to be somewhat tense. However, a minute later, he walks up to his teacher and hands her 80 cents. The teacher, amused, asks her what the extra 5 cents were for. The boy promptly replies, ""Teacher, this is a holy institution and there is no point in lying. While I was at it, I may have let one rip too."" ",A little boy in a very catholic school sharted and peed his pants...,0
post,3k41an,2qh72,jokes,false,1441730231,https://old.reddit.com/r/Jokes/comments/3k41an/sex_if_like_a_box_of_chocolate/,self.jokes,,You gotta check underneath to see what you're going to get.,Sex if like a box of chocolate...,0
post,3k40vp,2qh72,jokes,false,1441730061,https://old.reddit.com/r/Jokes/comments/3k40vp/whenever_somebody_hits_me_i_yell_somebody_grab/,self.jokes,,"""...I was just as**sa**u**lt**ed!""","Whenever somebody hits me, I yell, ""Somebody grab the pepper...""",0
post,3k3x94,2qh72,jokes,false,1441728571,https://old.reddit.com/r/Jokes/comments/3k3x94/my_friend_have_a_really_hot_mom_one_day_i_was/,self.jokes,,"Turns out his girlfriend is not answering his calls and he is on his way.
So I told his girlfriend turn on the phone and call him.",My friend have a really hot mom. One day I was having sex with his mom when he calls me and says he is on his way...,0
post,3k3wz8,2qh72,jokes,false,1441728457,https://old.reddit.com/r/Jokes/comments/3k3wz8/lpt_if_a_school_bully_is_tormenting_you_just/,self.jokes,,...otherwise he might spit in your burger later on in life.,"LPT: If a school bully is tormenting you, just ignore him...",1
post,3k3uh0,2qh72,jokes,false,1441727423,https://old.reddit.com/r/Jokes/comments/3k3uh0/how_many_redditors_does_it_take_to_screw_in_a_new/,self.jokes,,Zero. Somebody already did it.,How many redditors does it take to screw in a new lightbulb?,13
post,3k3ub8,2qh72,jokes,false,1441727360,https://old.reddit.com/r/Jokes/comments/3k3ub8/i_had_a_joke_about_insanity/,self.jokes,,but then I lost it.,I had a joke about insanity,12
post,3k3tx8,2qh72,jokes,false,1441727199,https://old.reddit.com/r/Jokes/comments/3k3tx8/i_hate_when_people_dont_finish_jokes/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k3tx8/i_hate_when_people_dont_finish_jokes/,,I hate when people don't finish jokes,0
post,3k3tbd,2qh72,jokes,false,1441726964,https://old.reddit.com/r/Jokes/comments/3k3tbd/an_officer_pulled_me_over_for_driving_erratically/,self.jokes,,He must have thought I was buzzed. ,"An officer pulled me over for driving erratically, but it was because some bees had gotten into my car.",8
post,3k3tas,2qh72,jokes,false,1441726958,https://old.reddit.com/r/Jokes/comments/3k3tas/did_you_know_that_youre_22_times_more_likely_to/,self.jokes,,[deleted],Did you know that you're 22 times more likely to be attacked by a cow than a shark?,5
post,3k3sza,2qh72,jokes,false,1441726827,https://old.reddit.com/r/Jokes/comments/3k3sza/why_us_didnt_attack_india_after_twintower/,self.jokes,,Because it didn't happen in 7/11,"Why US didn't attack India, after twin-tower incident, looking for terrorists ?",0
post,3k3suc,2qh72,jokes,false,1441726767,https://old.reddit.com/r/Jokes/comments/3k3suc/hey_guys_wanna_hear_a_joke/,self.jokes,,Reddit servers.,"Hey guys, wanna hear a joke?",3
post,3k3smw,2qh72,jokes,false,1441726653,https://old.reddit.com/r/Jokes/comments/3k3smw/i_got_catcalled_by_the_garbagemen_outside_my/,self.jokes,,They know a good piece of trash when they see one.  ,I got catcalled by the garbagemen outside my house this morning...,14
post,3k3s1b,2qh72,jokes,false,1441726415,https://old.reddit.com/r/Jokes/comments/3k3s1b/two_tomatoes_are_sitting_in_a_refrigerator/,self.jokes,,"One turns to the other and says: ""It's really cold in here"".

and the other one says:

[""JESUS CHRIST A TALKING TOMATO!!""](/spoiler)",Two tomatoes are sitting in a refrigerator,1
post,3k3r01,2qh72,jokes,false,1441725996,https://old.reddit.com/r/Jokes/comments/3k3r01/so_the_bass_clef_said_to_the_treble_clef/,self.jokes,,Don't take that tone with me,So the bass clef said to the treble clef,31
post,3k3qgz,2qh72,jokes,false,1441725777,https://old.reddit.com/r/Jokes/comments/3k3qgz/the_husband_comes_back_late_home_wife_greets_him/,self.jokes,," ""Where were you all this time?"", She asks him.
""I was playing chess with Tom"".
""And why do you smell of alcohol??"" she asks again, angrily.
husband replies "" What do you want me to smell like, chess?""
",The husband comes back late home... Wife greets him at the door..,0
post,3k3qg4,2qh72,jokes,false,1441725769,https://old.reddit.com/r/Jokes/comments/3k3qg4/my_wife_just_asked_me_what_i_think_about_syria/,self.jokes,,"I replied: ""Well, apart from Juventus or Roma I can't really see anyone else winning it this season""",My wife just asked me what I think about Syria,4
post,3k3qd7,2qh72,jokes,false,1441725728,https://old.reddit.com/r/Jokes/comments/3k3qd7/ten_dollars_is_ten_dollars/,self.jokes,,"Stumpy and his wife Martha went to the state fair every year. Every year Stumpy would say, ""Martha, I'd like to ride in that there airplane.""
And every year Martha would say, ""I know Stumpy, but that airplane ride costs ten dollars, and ten dollars is ten dollars.""


One year Stumpy and Martha went to the fair and Stumpy said, ""Martha, I'm 71 years old. If I don't ride that airplane this year I may never get another chance.""
Martha replied, ""Stumpy, that there airplane ride costs ten dollars, and ten dollars is ten dollars.""
The pilot overheard them and said, ""Folks, I'll make you a deal, I'll take you both up for a ride. If you can stay quiet for the entire ride and not say one word, I won't charge you, but if you say one word it's ten dollars.""
Stumpy and Martha agreed and up they went.


The pilot did all kinds of twists and turns, rolls and dives, but not a word was heard.
He did all his tricks over again, but still not a word.
They landed and the pilot turned to Stumpy, ""By golly, I did everything I could think of to get you to yell out, but you didn't."" Stumpy replied, ""Well, I was gonna say something when Martha fell out, but ten dollars is ten dollars."" 

edit--format",Ten dollars is ten dollars.,3893
post,3k3pr5,2qh72,jokes,false,1441725466,https://old.reddit.com/r/Jokes/comments/3k3pr5/til_a_study_revealed_that_users_never_check_the/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k3pr5/til_a_study_revealed_that_users_never_check_the/,,TIL: A study revealed that users never check the authenticity of facts they find on /r/todayilearned,3
post,3k3pq0,2qh72,jokes,false,1441725450,https://old.reddit.com/r/Jokes/comments/3k3pq0/how_do_you_keep_an_idiot_in_suspense_for_24_hours/,self.jokes,,I'll tell you the answer tomorrow.,How do you keep an idiot in suspense for 24 hours?,1
post,3k3poc,2qh72,jokes,false,1441725429,https://old.reddit.com/r/Jokes/comments/3k3poc/a_man_was_afraid_to_go_into_kohls_at_the_local/,self.jokes,,"because according to the sign:

Kohls

Staples

Dicks",A man was afraid to go into Kohl's at the local strip mall,0
post,3k3pec,2qh72,jokes,false,1441725308,https://old.reddit.com/r/Jokes/comments/3k3pec/my_girlfriend_treats_me_like_a_god/,self.jokes,,She takes little notice of my existence unless she wants something.,My girlfriend treats me like a God,233
post,3k3p9k,2qh72,jokes,false,1441725251,https://old.reddit.com/r/Jokes/comments/3k3p9k/about_the_newest_microsoft_patch/,self.jokes,,"Microsoft confirms that there's an issue with their most recent patch: it can corrupt Windows installations.  A Microsoft developer by the name of Benedict [Last name withheld due to reddit rules] admitted that the code he wrote was faulty and could lead to corruption of some system files.   
However, Microsoft still recommends downloading the patch, since these cases are rare, and a tool that repairs affected installations will be available by tomorrow, and can easily be downloaded, since the faulty patch doesn't break any Internet features.  Microsoft estimates that only 0.002% of Windows installations will be affected, and that on all other PCs, the patch does fix the bug it addresses.  Although some sources on the net claim otherwise, Microsoft states that...

Benedict's Blunder Patch is low-key.",About the newest Microsoft patch,1
post,3k3o8w,2qh72,jokes,false,1441724819,https://old.reddit.com/r/Jokes/comments/3k3o8w/prematurely_born/,self.jokes,,[deleted],Prematurely born.,0
post,3k3o25,2qh72,jokes,false,1441724737,https://old.reddit.com/r/Jokes/comments/3k3o25/have_you_ever_spelt_a_hard_word_with_so_much/,self.jokes,,[deleted],Have you ever spelt a hard word with so much confidence that even auto correct took a extra minute to realize it was spelt wrong.,0
post,3k3non,2qh72,jokes,false,1441724586,https://old.reddit.com/r/Jokes/comments/3k3non/a_kindergarten_teacher_asks_her_students_what/,self.jokes,,"She said, ""What does a chicken give us?"" and the students replied, ""Eggs"". She then asked, ""What does a pig give us?"" and the students replied a joyous ""Bacon"". Finally she asked ""What does a cow give us?"" and before anyone could answer little Johnny said ""Homework"".

Joke provided by my ten year old son.",A kindergarten teacher asks her students what animals provide us...,249
post,3k3nhd,2qh72,jokes,false,1441724496,https://old.reddit.com/r/Jokes/comments/3k3nhd/i_tried_to_give_my_cat_a_bath/,self.jokes,,[deleted],I tried to give my cat a bath...,7
post,3k3mns,2qh72,jokes,false,1441724138,https://old.reddit.com/r/Jokes/comments/3k3mns/in_america_child_protection_saves_your_kids_from/,self.jokes,,In Soviet Russia child protection beats your kids ,In America child protection saves your kids from your beating,0
post,3k3m9i,2qh72,jokes,false,1441723973,https://old.reddit.com/r/Jokes/comments/3k3m9i/reddit_servers/,self.jokes,,[deleted],Reddit Servers.,2
post,3k3l76,2qh72,jokes,false,1441723414,https://old.reddit.com/r/Jokes/comments/3k3l76/the_dirtiest_one_of_them_all/,self.jokes,,A pale white horse galloped and jumped into muddy water,The dirtiest one of them all,0
post,3k3l5l,2qh72,jokes,false,1441723397,https://old.reddit.com/r/Jokes/comments/3k3l5l/are_you_a_democrat_republican_or_a_southerner/,self.jokes,,"Are you a Democrat, Republican, or a Southerner?  Here is a little test that will help you decide.  The answer can be found by posing the following question:

*You’re walking down the street with your husband/wife and your two small children.  Suddenly, an Islamic Terrorist with a huge knife comes around the corner, locks eyes with you, screams obscenities, praises Allah, raises the
knife, and charges at you. You are carrying a Glock 40 caliber. What do you do?*


**The Democrat’s Answer:**

Well, that’s not enough information to answer the question!
Does the man look poor or oppressed?
Have I ever done anything to him that would inspire him to attack?
Could we run away?
What does my wife/husband think?
What about the kids?
Could I possibly swing the gun like a club and knock the knife out of his hand?
What does the law say about this situation?
Does the Glock have appropriate safety built into it?
Why am I carrying a loaded gun anyway, and what kind of message does this send to society and to my children?
Is it possible he’d be happy with just killing me?
Does he definitely want to kill me, or would he be content just to wound me?
If I were to grab his knees and hold on, could my family get away while he was stabbing me?
Should I call 9-1-1?
Why is this street so deserted?
We need to raise taxes, have a paint and weed day, and make this happier, healthier street that would discourage such behavior.
This is all so confusing! I need to debate this with some friends for few days and try to come to a consensus.

**The Republican’s Answer:**

BANG!


**The Southerner’s Answer:**

BANG! BANG! BANG! BANG! BANG! BANG! BANG! BANG!

BANG! Click….. (Sounds of reloading)

BANG! BANG! BANG!

BANG! BANG! BANG! BANG! BANG!

BANG! Click

Daughter: “Nice grouping, Daddy! Were those the Winchester Silver Tips or
Hollow Points?”

Son: “Can I shoot the next one!??!”

Wife: “You ain’t taking that to the Taxidermist!”","Are you a Democrat, Republican or a Southerner?",3
post,3k3kwv,2qh72,jokes,false,1441723292,https://old.reddit.com/r/Jokes/comments/3k3kwv/once_upon_a_timethere_was_this_cute_black_rabbit/,self.jokes,,...he used to breath from his arsehole.After a long day of collecting carrots he sat down to rest and died.,"Once upon a time,there was this cute black rabbit...",0
post,3k3kdp,2qh72,jokes,false,1441723064,https://old.reddit.com/r/Jokes/comments/3k3kdp/i_was_arrested_for_shoplifting_the_other_day/,self.jokes,,"I had to explain to the officer that it was all a misunderstanding, I was attempting to pick up the eggs which were free, I just don't know what ""range eggs"" are.",I was arrested for shoplifting the other day,0
post,3k3k9z,2qh72,jokes,false,1441723011,https://old.reddit.com/r/Jokes/comments/3k3k9z/the_blind_pilots/,self.jokes,,"Passengers of a 747 begin settling in for their scheduled takeoff when two men in pilot uniforms stumble into the plane, one with a seeing eye dog and the other with a walking stick.  The passengers think it's some sort of joke and think nothing of it, but the men carefully and methodically make their way to the cockpit.

The passengers look at each other a little uneasy but say nothing.  The plane starts down the runway ever-increasing in speed.  The passengers see the end of the runway approaching and start to mumble to themselves.  The plane doesn't pull up and the runaway end comes ever nearer.  A couple passengers release muffled screams and begin to panic, but the plane continues to the end of the runaway.  The passengers at this point begin a full-blown panic and scream loudly and right before they hit the trees at the end of the runway, the plane lifts off without a hitch just barely grazing the tops of the trees as it passes.

Inside the cockpit, the blind copilot turns to the other and says, ""That was close.  You know one day they're not gonna scream and we're all gonna die.""",The blind pilots,680
post,3k3k7i,2qh72,jokes,false,1441722984,https://old.reddit.com/r/Jokes/comments/3k3k7i/what_vocation_can_transform_anything_into_a_gate/,self.jokes,,A reporter.,What vocation can transform anything into a gate?,1
post,3k3juh,2qh72,jokes,false,1441722829,https://old.reddit.com/r/Jokes/comments/3k3juh/8_shot_mag/,self.jokes,,"A guy walked  into a crowded bar, waving his UN-holstered pistol and  yelled,  I have a .45 Colt with an eight-shot magazine and  I want to know who's been sleeping with my wife.""
 
A voice from the back of the room called out,   You don't have enough ammo!""
",8 shot mag,1
post,3k3jik,2qh72,jokes,false,1441722689,https://old.reddit.com/r/Jokes/comments/3k3jik/opinions_are_like_assholes/,self.jokes,,[deleted],Opinions are like assholes...,1
post,3k3jhd,2qh72,jokes,false,1441722678,https://old.reddit.com/r/Jokes/comments/3k3jhd/a_man_was_driving_down_the_road/,self.jokes,,[deleted],A man was driving down the road...,51
post,3k3i4q,2qh72,jokes,false,1441722096,https://old.reddit.com/r/Jokes/comments/3k3i4q/i_was_driving_recklessly_around_the_city_and/,self.jokes,,"She said, ""Hey! You wanna smash me?""

I said, ""Sorry babe. Don't have a condom right now, maybe later.""",I was driving recklessly around the city and almost hit a hot girl,0
post,3k3hgs,2qh72,jokes,false,1441721810,https://old.reddit.com/r/Jokes/comments/3k3hgs/why_did_the_skeletons_start_dancing/,self.jokes,,Because they forgot the g in graveyard.,Why did the skeletons start dancing?,0
post,3k3gxm,2qh72,jokes,false,1441721590,https://old.reddit.com/r/Jokes/comments/3k3gxm/how_do_chemists_get_high/,self.jokes,,they drop acid of course,How do chemists get high?,0
post,3k3gje,2qh72,jokes,false,1441721405,https://old.reddit.com/r/Jokes/comments/3k3gje/what_would_people_call_an_old_john_cena/,self.jokes,,John Senile,What would people call an old John Cena?,0
post,3k3g7y,2qh72,jokes,false,1441721258,https://old.reddit.com/r/Jokes/comments/3k3g7y/so_we_were_having_a_religious_appreciation_day_in/,self.jokes,,"The professor says ""if you're Catholic please stand!"" 

a few people stand

The professor says ""Baptist please stand"" 

Going to school in the south of course the majority stands 

The professor says ""If you're Jewish please stand."" 

And I yell, ""We're not falling for that again!"" 

I know it's not too funny but I hope it made ya smile a bit",So we were having a religious appreciation day in class today,13
post,3k3g11,2qh72,jokes,false,1441721158,https://old.reddit.com/r/Jokes/comments/3k3g11/ever_wonder_why_tiny_little_paper_cuts_hurt_so_bad/,self.jokes,,Cause you're a pussy,Ever wonder why tiny little paper cuts hurt so bad?,1
post,3k3ee3,2qh72,jokes,false,1441720407,https://old.reddit.com/r/Jokes/comments/3k3ee3/why_was_6_afraid_of_7/,self.jokes,,[deleted],Why was 6 afraid of 7?,0
post,3k3eda,2qh72,jokes,false,1441720400,https://old.reddit.com/r/Jokes/comments/3k3eda/i_got_kicked_out_of_the_chorus_line_i_was_with/,self.jokes,,I just couldn’t stay in sequins.,I got kicked out of the chorus line I was with.,0
post,3k3dyc,2qh72,jokes,false,1441720190,https://old.reddit.com/r/Jokes/comments/3k3dyc/우리카지노ask237com쿠폰확실하게챙겨드립니다/,self.jokes,,[removed],우리카지노&lt;Ask237.com&gt;&lt;쿠폰확실하게챙겨드립니다&gt;,1
post,3k3bln,2qh72,jokes,false,1441719030,https://old.reddit.com/r/Jokes/comments/3k3bln/shot_my_first_turkey_today/,self.jokes,,Scared everyone in the frozen meat department. ,Shot my first turkey today.,80
post,3k3b4q,2qh72,jokes,false,1441718806,https://old.reddit.com/r/Jokes/comments/3k3b4q/what_did_the_astronaut_say_to_his_girlfriend_when/,self.jokes,,I need some space.,What did the astronaut say to his girlfriend when he broke up with her?,33
post,3k3amc,2qh72,jokes,false,1441718590,https://old.reddit.com/r/Jokes/comments/3k3amc/in_light_of_germanys_discovery_of_isis_using/,self.jokes,,"What do you call a soldier who's survived mustard gas and pepper spray? 

A seasoned veteran.",In light of Germany's discovery of ISIS using mustard gas:,9
post,3k39r1,2qh72,jokes,false,1441718190,https://old.reddit.com/r/Jokes/comments/3k39r1/i_was_walking_down_the_street_one_day_and_stepped/,self.jokes,,[deleted],I was walking down the street one day and stepped on something soft...,1
post,3k390z,2qh72,jokes,false,1441717744,https://old.reddit.com/r/Jokes/comments/3k390z/what_is_the_biggest_crime_committed_by/,self.jokes,,Male fraud.,What is the biggest crime committed by transvestites?,21
post,3k38hh,2qh72,jokes,false,1441717473,https://old.reddit.com/r/Jokes/comments/3k38hh/war_is_gods_way_of_teaching_americans_geography/,self.jokes,,[deleted],War is God's way of teaching Americans geography.,1
post,3k38ez,2qh72,jokes,false,1441717440,https://old.reddit.com/r/Jokes/comments/3k38ez/what_drink_does_hitler_hate_the_most/,self.jokes,,Juice,What drink does hitler hate the most?,2
post,3k388s,2qh72,jokes,false,1441717360,https://old.reddit.com/r/Jokes/comments/3k388s/whats_the_difference_between_a_gay_man_a/,self.jokes,,[deleted],Whats the difference between a gay man &amp; a refrigerator?,4
post,3k384m,2qh72,jokes,false,1441717304,https://old.reddit.com/r/Jokes/comments/3k384m/did_you_hear_about_the_guy_who_used_to_date_a/,self.jokes,,[deleted],Did you hear about the guy who used to date a pizza?,0
post,3k383r,2qh72,jokes,false,1441717290,https://old.reddit.com/r/Jokes/comments/3k383r/rape_game/,self.jokes,,"Husband: Darling, let's play rape game

Wife: No!

Husband: Perfect start ",Rape game,1
post,3k3783,2qh72,jokes,false,1441716655,https://old.reddit.com/r/Jokes/comments/3k3783/before_it_starts/,self.jokes,,"
A man comes home from an exhausting day at work, plops down on the couch in front of the television, and tells his wife, ""Get me a beer before it starts."" The wife sighs and gets him a beer. Fifteen minutes later, the man says, ""Get me another beer before it starts."" She looks cross, but fetches another beer and slams it down next to him. He finishes that beer and a few minutes later says, ""Quick, get me another beer, it's going to start any minute."" The wife is furious. She yells at him, ""Is that all you're going to do tonight? Drink beer and sit in front of that TV? You’re nothing but a lazy, drunken, fat slob."" The man sighs and says, ""It’s started…""
",BEFORE IT STARTS,238
post,3k36on,2qh72,jokes,false,1441716369,https://old.reddit.com/r/Jokes/comments/3k36on/what_do_you_take_to_an_ethiopian_wedding/,self.jokes,,[deleted],What do you take to an Ethiopian wedding?,0
post,3k36ff,2qh72,jokes,false,1441716243,https://old.reddit.com/r/Jokes/comments/3k36ff/whats_the_difference_between_a_bdsm_slavegirl_and/,self.jokes,,The mosquito stops sucking if you slap it. ,"Whats the difference between a bdsm slavegirl, and a mosquito?",108
post,3k36cq,2qh72,jokes,false,1441716205,https://old.reddit.com/r/Jokes/comments/3k36cq/as_football_starts_id_just_like_to_give_players_a/,self.jokes,,[deleted],"As football starts , I'd just like to give players a tip.",4
post,3k36ce,2qh72,jokes,false,1441716200,https://old.reddit.com/r/Jokes/comments/3k36ce/jamaican_space_program/,self.jokes,,Have you heard of the Jamaican space program? they just keep getting higher and higher and higher......,Jamaican space program.,2
post,3k369t,2qh72,jokes,false,1441716171,https://old.reddit.com/r/Jokes/comments/3k369t/i_told_my_friends_i_had_a_date_with_a_really/,self.jokes,,[deleted],I told my friends I had a date with a really attractive girl,0
post,3k3639,2qh72,jokes,false,1441716078,https://old.reddit.com/r/Jokes/comments/3k3639/an_irshman_leaves_a_bar/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k3639/an_irshman_leaves_a_bar/,,An Irshman leaves a bar.,11
post,3k34k5,2qh72,jokes,false,1441715167,https://old.reddit.com/r/Jokes/comments/3k34k5/jokes/,self.jokes,,[removed],JOKES,1
post,3k34bg,2qh72,jokes,false,1441715036,https://old.reddit.com/r/Jokes/comments/3k34bg/a_guy_and_his_wife_are_sitting_and_watching_a/,self.jokes,,[deleted],A guy and his wife are sitting and watching a boxing match on television.,0
post,3k33pi,2qh72,jokes,false,1441714712,https://old.reddit.com/r/Jokes/comments/3k33pi/two_alligators_in_dc/,self.jokes,,[deleted],Two Alligators in DC,0
post,3k322r,2qh72,jokes,false,1441713749,https://old.reddit.com/r/Jokes/comments/3k322r/who_let_the_docs_out/,self.jokes,,Google. Google docs.,Who let the docs out?,0
post,3k2zxl,2qh72,jokes,false,1441712384,https://old.reddit.com/r/Jokes/comments/3k2zxl/why_did_the_chicken_cross_the_road/,self.jokes,,[deleted],^Why did the chicken cross the road?,1
post,3k2zgc,2qh72,jokes,false,1441712077,https://old.reddit.com/r/Jokes/comments/3k2zgc/lost_my_watch_at_a_party/,self.jokes,,[deleted],Lost my watch at a party...,0
post,3k2xuy,2qh72,jokes,false,1441710972,https://old.reddit.com/r/Jokes/comments/3k2xuy/if_you_dont_drink/,self.jokes,,"...then all of your stories suck and end with, ""And then I got home""",If you don't drink...,0
post,3k2xtj,2qh72,jokes,false,1441710948,https://old.reddit.com/r/Jokes/comments/3k2xtj/if_panic_at_the_disco_were_mexican/,self.jokes,,They would be called Hispanics at the disco,If Panic! At the disco were Mexican...,2
post,3k2xlk,2qh72,jokes,false,1441710800,https://old.reddit.com/r/Jokes/comments/3k2xlk/during_loving_father_to_mom_i_said_dont_and_got/,self.jokes,,[removed],"During loving father to mom, i said don't and got reply who are you?",1
post,3k2xlb,2qh72,jokes,false,1441710793,https://old.reddit.com/r/Jokes/comments/3k2xlb/im_planning_a_marriage_proposal_over_the_phone/,self.jokes,,[deleted],I'm planning a marriage proposal over the phone.,3
post,3k2xd1,2qh72,jokes,false,1441710640,https://old.reddit.com/r/Jokes/comments/3k2xd1/ahh_mexico/,self.jokes,,The silver metal winner of the Mexican-American War.,Ahh Mexico...,0
post,3k2wt3,2qh72,jokes,false,1441710282,https://old.reddit.com/r/Jokes/comments/3k2wt3/asdasd/,self.jokes,,[removed],asdasd,0
post,3k2wgk,2qh72,jokes,false,1441710058,https://old.reddit.com/r/Jokes/comments/3k2wgk/what_did_the_police_officer_say_to_the_iphone_who/,self.jokes,,You are charged with Battery,What did the police officer say to the iPhone who abused his wife?,0
post,3k2w9c,2qh72,jokes,false,1441709926,https://old.reddit.com/r/Jokes/comments/3k2w9c/i_decided_to_put_some_ketchup_in_my_eyes/,self.jokes,,"...but in Heinzsight, it wasn't a good idea.",I decided to put some ketchup in my eyes...,73
post,3k2vw8,2qh72,jokes,false,1441709656,https://old.reddit.com/r/Jokes/comments/3k2vw8/man_goes_to_the_doctor/,self.jokes,,"""Doc, doc, the area around the entrance on my butt is a little itchy""

""I think you mean the exit.........""",Man goes to the doctor,0
post,3k2vuc,2qh72,jokes,false,1441709621,https://old.reddit.com/r/Jokes/comments/3k2vuc/imgbbnet_earn_up_to_61000_views_paypal_btc/,self.jokes,,[removed],"ImgBB.net - Earn up to 6$/1000 views - Paypal, BTC, Payonner, Payza, Skrill, WMZ",1
post,3k2vu3,2qh72,jokes,false,1441709614,https://old.reddit.com/r/Jokes/comments/3k2vu3/my_friend_met_daniel_craig_at_a_bar_last_night_he/,self.jokes,,She said it was decent Bondage.,"My friend met Daniel Craig at a bar last night. He took her back to his, handcuffed her, tied her to the bedposts and fucked her brains out...",0
post,3k2usr,2qh72,jokes,false,1441708876,https://old.reddit.com/r/Jokes/comments/3k2usr/things_south_africans_do/,self.jokes,,"You’re working on your computer and you’re in the habit of clicking ‘SAVE’ very often, in case of load shedding

You speed up for an orange robot, not traffic light

You check the robots before you go when they turn green in case a taxi is still going through red

Travelling at 120 km/h, you’re the slowest vehicle on the freeway

The first thing you do when you get in your car is lock the doors

You produce a R100 note instead of your driver’s licence when stopped by a traffic officer

You flash your brights at oncoming traffic to warn them about a speed cop trapping in the bushes

You prefer private transport to public transport, because taking a taxi means sharing a lift with 40 people

You love the fact that we have 11 official languages, even though you can only speak one or two of them



You can sing your national anthem in four languages and you have no idea what it means in any of them

Some of your fellow citizens have the most festive names, such as Blessing, Christmas, Innocence, Precious, Gift, Patience, Pretty

You don’t say ‘yes’, you say ‘ja’ or ‘yebo’

You always say ‘ja no definitely’

You put ‘man’ at the end of every sentence

You SMS your chommie, not text (well now you WhatsApp)

You’ve had at least one thing stolen from you

You love how Zapiro always gets it right

You have an opinion about the Oscar Pistorius case",Things South Africans Do…,0
post,3k2tch,2qh72,jokes,false,1441707817,https://old.reddit.com/r/Jokes/comments/3k2tch/what_do_you_call_a_biscuit_on_a_motorbike/,self.jokes,,A bikkie.,What do you call a biscuit on a motorbike?,0
post,3k2sr8,2qh72,jokes,false,1441707377,https://old.reddit.com/r/Jokes/comments/3k2sr8/you_can_tell_the_gender_of_an_ant_by_putting_it/,self.jokes,,"If it sinks: Girl Ant


If it floats: Boy ant",You can tell the gender of an Ant by putting it in water,22
post,3k2rkt,2qh72,jokes,false,1441706537,https://old.reddit.com/r/Jokes/comments/3k2rkt/why_is_it_once_you_go_black_you_never_go_back/,self.jokes,,Because no one will take you back ,Why is it once you go black you never go back?,0
post,3k2r37,2qh72,jokes,false,1441706180,https://old.reddit.com/r/Jokes/comments/3k2r37/what_time_did_the_star_trek_character_clone/,self.jokes,,[deleted],What time did the Star Trek character clone himself?,0
post,3k2oju,2qh72,jokes,false,1441704171,https://old.reddit.com/r/Jokes/comments/3k2oju/some_very_funny_adult_jokes/,self.jokes,,[removed],Some Very Funny Adult Jokes !!!,1
post,3k2nkj,2qh72,jokes,false,1441703459,https://old.reddit.com/r/Jokes/comments/3k2nkj/in_a_room_of_engineers_how_many_does_it_take_to/,self.jokes,,"All of them.

However, it still hasn't been changed because they are each working on a more efficient bulb and thread, followed by a lot of arguing.","In a room of engineers, how many does it take to screw in a light bulb?",0
post,3k2mza,2qh72,jokes,false,1441703029,https://old.reddit.com/r/Jokes/comments/3k2mza/whats_the_best_thing_about_having_insomnia/,self.jokes,,Only one nights sleep til Christmas!,What's the best thing about having insomnia?,22
post,3k2mpd,2qh72,jokes,false,1441702841,https://old.reddit.com/r/Jokes/comments/3k2mpd/has_this_been_posted_before/,self.jokes,,Has this been posted before?,Has this been posted before?,0
post,3k2mfp,2qh72,jokes,false,1441702641,https://old.reddit.com/r/Jokes/comments/3k2mfp/why_the_chicken_crossed_the_road/,self.jokes,,"RONALD FISHER: Why does it have to be a chicken? Why not a frog, turkey, or pig? We randomly try to a have chicken, frog, turkey and pig cross the road 10 times each. We then compare the mean number of times each animal crossed the road to determine if there's a difference in means. 

SARAH PALIN: The chicken crossed the road because, gosh-darn it, he's a maverick!

BARACK OBAMA: The chicken crossed the road because it was time for change! The chicken wanted change! 

JOHN McCAIN: My friends, that chicken crossed the road because he recognized the need to engage in cooperation and dialogue with all the chickens on the other side of the road.

HILLARY CLINTON: When I was First Lady, I personally helped that little chicken to cross the road. This experience makes me uniquely qualified to ensure right from Day One that every chicken in this country gets the chance it deserves to cross the road. But then, this really isn't about me.

GEORGE W. BUSH: We don't really care why the chicken crossed the road. We just want to know if the chicken is on our side of the road, or not. The chicken is either against us, or for us. There is no middle ground here.

DICK CHENEY: Where's my gun?

COLIN POWELL: Now to the left of the screen, you can clearly see the satellite image of the chicken crossing the road. 

BILL CLINTON: I did not cross the road with that chicken. 

JOHN KERRY: Although I voted to let the chicken cross the road, I am now against it! It was the wrong road to cross, and I was misled about the chicken's intentions. I am not for it now, and will remain against it. 

DR. PHIL: The problem we have here is that this chicken won't realize that he must first deal with the problem on this side of the road before it goes after the problem on the other side of the road. What we need to do is help him realize how stupid he's acting by not taking on his current problems before adding new problems. 

OPRAH: Well, I understand that the chicken is having problems, which is why he wants to cross this road so bad. So instead of having the chicken learn from his mistakes and take falls, which is a part of life, I'm going to give this chicken a NEW CAR so that he can just drive across the road and not live his life like the rest of the chickens. 

NANCY GRACE: That chicken crossed the road because he's guilty! You can see it in his eyes and the way he walks. 

MARTHA STEWART: No one called me to warn me which way that chicken was going. I had a standing order at the Farmer's Market to sell my eggs when the price dropped to a certain level. No little bird gave me any insider information. 

JOHN LENNON: Imagine all the chickens in the world crossing roads together, in peace.

BILL GATES: I have just released eChicken2010, which will not only cross roads, but will lay eggs, file your important documents, and balance your checkbook. Internet Explorer is an integral part of eChicken2010. This new platform is much more stable and will never reboot. 

AUGUST MOBIUS: To get to the same side. 

ISAAC NEWTON: Chickens at rest tend to stay at rest. Chickens in motion tend to cross the road. 

WERNER HEISENBERG: We are not sure which side of the road the chicken was on, but it was moving very fast. 

DARTH VADER: Because it could not resist the power of the Dark Side. 

JERRY SEINFELD: Why does anyone cross a road? I mean, why doesn't anyone ever think to ask, ""What the heck was this chicken doing walking all over the place anyway?"" 

AL GORE: I will fight for the chickens and I will not disappoint them. Did I mention that I invented roads? 

KEN STARR: I intend to prove that the chicken crossed the road at the behest of the president of the United States of America in an effort to distract law enforcement officials and the American public from the criminal wrongdoing our highest elected official has been trying to cover up. As a result, the chicken is just another pawn in the president's ongoing and elaborate scheme to obstruct justice and undermine the rule of law. For that reason, my staff intends to offer the chicken unconditional immunity provided he cooperates fully with our investigation. Furthermore, the chicken will not be permitted to reach the other side of the road until our investigation and any Congressional follow-up investigations have been completed. 

PAT BUCHANAN: To steal a job from a decent, hardworking American. 

DR. SEUSS: Did the chicken cross the road? Did he cross it with a toad? Yes! The chicken crossed the road, but why it crossed, I've not been told! 

ERNEST HEMINGWAY: To die. In the rain. 

MARTIN LUTHER KING, JR.: I envision a world where all chickens will be free to cross roads without having their motives called into question. 

GRANDPA: In my day, we didn't ask why the chicken crossed the road. Someone told us that the chicken crossed the road, and that was good enough for us. 

ARISTOTLE: It is the nature of chickens to cross the road. 

KARL MARX: It was a historical inevitability. 

SADDAM HUSSEIN: This was an unprovoked act of rebellion and we were quite justified in dropping 50 tons of nerve gas on it. 

RONALD REAGAN: What chicken? 

CAPTAIN JAMES T. KIRK: To boldly go where no chicken has gone before. 
FOX MULDER: You saw it cross the road with your own eyes. How many more chickens have to cross before you believe it? 

MACHIAVELLI: The point is that the chicken crossed the road. Who cares why? The end of crossing the road justifies whatever motive there was. 
FREUD: The fact that you are at all concerned that the chicken crossed the road reveals your underlying sexual insecurity. 

ALBERT EINSTEIN: Did the chicken really cross the road or did the road move beneath the chicken? 

IMMANUEL KANT: The chicken was acting out of a sense of duty to cross the road, as chickens have traditionally crossed roads throughout history. 

THE BIBLE: And God came down from the heavens, and He said unto the chicken, ""Thou shalt cross the road."" And the chicken crossed the road, and there was much rejoicing. 

COLONEL SANDERS: I missed one? 
RICHARD M. NIXON: The chicken did not cross the road. I repeat, the chicken did not cross the road. I don't know any chickens. I have never known any chickens. 

JANOS von NEUMANN: The chicken is distributed probabilistically on all sides of the road until you observe it on your side. 

BARBARA WALTERS: Isn't that interesting? In a few moments, we will be listening to the chicken tell, for the first time, the heart warming story of how it experienced a serious case of molting, and went on to accomplish its life long dream of crossing the road. 

ANDERSON COOPER, CNN: We have reason to believe there is a chicken, but we have not yet been allowed to have access to the other side of the road. 

DONALD RUMSFELD: Now to the left of the screen, you can clearly see the satellite image of the chicken crossing the road. 

ANDRE AMPERE: To keep up with current events. 

ROBERT BOYLE: She had been under too much pressure at home. 

JAMES WATT: It thought it would be a good way to let off steam. 

THOMAS EDISON: She thought it would be an illuminating experience. 

JEAN FOUCALT: It didn't. The rotation of the earth made it appear to cross. 
KARL GAUSS: Because of the magnetic personality of the rooster on the other side. 

GUSATV HERTZ: Lately, its been crossing with greater frequency. 

GEORG OHM: There was more resistance on this side of the road. 

ERWIN SCHRODINGER: Since the wording of the question implies the absence of an observer (else the fowl's motivation might easily be deduced), it is evident that the chicken simultaneously did and did not cross the road. In the face of this, any speculation as to the bird's purpose must be viewed as mere sophistry - and as such is beyond the bounds of this discussion.",Why the chicken crossed the road,3
post,3k2m1b,2qh72,jokes,false,1441702285,https://old.reddit.com/r/Jokes/comments/3k2m1b/how_do_you_know_the_passengers_of_the_missing/,self.jokes,,A new season of lost is out now!,How do you know the passengers of the missing plane are alive?,0
post,3k2lzz,2qh72,jokes,false,1441702258,https://old.reddit.com/r/Jokes/comments/3k2lzz/putin_goes_on_holiday/,self.jokes,,"Vladimir Putin arrives at an airport, gets in line at customs desk.
Customs officer: Occupation?
Putin: No, just visiting.",Putin goes on holiday!,26
post,3k2kuf,2qh72,jokes,false,1441701324,https://old.reddit.com/r/Jokes/comments/3k2kuf/i_accidentally_bought_a_bicycle_that_has_no_seat/,self.jokes,,it's not a deal breaker but it's kind of a pain in the ass.,I accidentally bought a bicycle that has no seat,14
post,3k2iz2,2qh72,jokes,false,1441699794,https://old.reddit.com/r/Jokes/comments/3k2iz2/one_man_gave_his_life_so_you_could_have/,self.jokes,,🎺 🎺 🎺 🎺 JOHN CENA 🎺 🎺 🎺 🎺,"One man gave his life, so you could have everything you ever wanted, and his name was",0
post,3k2iz0,2qh72,jokes,false,1441699793,https://old.reddit.com/r/Jokes/comments/3k2iz0/hillary_and_mandela/,self.jokes,,"Poor Hillary was down in the dumps this morning, the campaign is in the doldrums, the pollsters are not being kind, the public is disinterested, and she is way behind in New Hampshire. To top it all off, now she is even having to consider Joe Biden as a potential competitor. Uncle Joe Biden! For crying out loud.




So Bill did his best to try to cheer her up this morning, over breakfast. He reminded her of their good acquaintance, Nelson Mandela, who faced even greater hardship and adversities in his life, but still overcame them and triumphed. And he reminded her to look on the bright side: Nelson Mandela was elected President after he was released from prison.",Hillary and Mandela,1
post,3k2i1e,2qh72,jokes,false,1441699135,https://old.reddit.com/r/Jokes/comments/3k2i1e/what_does_a_gas_discharge_lamp/,self.jokes,,Fart fart fart XD,What does a gas discharge lamp?,0
post,3k2i0a,2qh72,jokes,false,1441699104,https://old.reddit.com/r/Jokes/comments/3k2i0a/bruce_willis/,self.jokes,,"Bruce Willis will probably keep making action movies. Because, you know what they say about old habits...",Bruce Willis...,1
post,3k2hpk,2qh72,jokes,false,1441698851,https://old.reddit.com/r/Jokes/comments/3k2hpk/what_do_you_call_blackman_in_disguise/,self.jokes,,[deleted],What do you call blackman in disguise?,0
post,3k2h7v,2qh72,jokes,false,1441698480,https://old.reddit.com/r/Jokes/comments/3k2h7v/everybody_keeps_downvoting_my_racist_jokes/,self.jokes,,It's like a load of black people have suddenly gotten laptops or something.,Everybody keeps downvoting my racist jokes,0
post,3k2g72,2qh72,jokes,false,1441697679,https://old.reddit.com/r/Jokes/comments/3k2g72/what_does_a_light_bulb_filled_with_gas/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k2g72/what_does_a_light_bulb_filled_with_gas/,,What does a light bulb filled with gas?,0
post,3k2f7i,2qh72,jokes,false,1441696903,https://old.reddit.com/r/Jokes/comments/3k2f7i/if_terminator_had_a_horse_what_would_its_name_be/,self.jokes,,"Termineightor



I'll show myself out...","If Terminator had a horse, what would its name be?",3
post,3k2eiq,2qh72,jokes,false,1441696415,https://old.reddit.com/r/Jokes/comments/3k2eiq/what_do_you_call_someone_without_a_nose_or_a_body/,self.jokes,,"Nobody nose.

Source: Anonymous",What do you call someone without a nose or a body?,5
post,3k2ehe,2qh72,jokes,false,1441696388,https://old.reddit.com/r/Jokes/comments/3k2ehe/joke_what_does_a_light_bulb_filled_with_gas/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k2ehe/joke_what_does_a_light_bulb_filled_with_gas/,,(JOKE) What does a light bulb filled with gas?,0
post,3k2d15,2qh72,jokes,false,1441695380,https://old.reddit.com/r/Jokes/comments/3k2d15/til_that_it_is_estimated_that_up_to_90_of_people/,self.jokes,,[deleted],TIL that it is estimated that up to 90% of people in the US will begin to read a post without checking the subreddit it's posted in.,1
post,3k2cpb,2qh72,jokes,false,1441695126,https://old.reddit.com/r/Jokes/comments/3k2cpb/what_do_you_tell_a_cow_thats_in_the_way/,self.jokes,,Mooooooooooooove. ,What do you tell a cow that's in the way?,0
post,3k2c26,2qh72,jokes,false,1441694687,https://old.reddit.com/r/Jokes/comments/3k2c26/why_is_sia_not_in_her_music_videos/,self.jokes,,Because she doesn't want anyone to Sia,Why is Sia not in her music videos?,6
post,3k2aj5,2qh72,jokes,false,1441693585,https://old.reddit.com/r/Jokes/comments/3k2aj5/i_just_found_out_that_the_reptile_i_had_sex_with/,self.jokes,,Now I have a dino-sore,I just found out that the reptile I had sex with last night had an STD,0
post,3k29cd,2qh72,jokes,false,1441692749,https://old.reddit.com/r/Jokes/comments/3k29cd/3_nuns_are_at_the_pearly_gates/,self.jokes,,"St Peter greets them saying ""Sisters of the faith! I have some bad news. Due to the current state of the world, there is a lineup to get into heaven. But since you devoted your lives to the Lord, I have a special surprise for you! You all get to go back to Earth until we can get you in past the gates! And the best part is, because you lived a life of sacrifice and poverty, we will let you return as any famous or rich person you want! Isn't that great?!""

He looks to the first nun, ""Who would you like to be?""
""I want to be Madonna, in 1987. She could really dance!""
POOF! She is sent down below.

""And you?"" St. Peter says, looking at the second nun.
""I want to be Oprah. She has a good heart, and more money than I can spend I'm sure!""
POOF! She's on her way.

""And you?"" he says, looking at the final nun.
In her thick Italian accent, she struggles with the words, ""Alberto Peepalini""

St Peter looks confused, and begins to search through his scrolls. Nowhere does he find this Alberto character. ""Sister, are you sure you have the name right? I can't find a record of him...""

""Yes! I can prove it!"" she says, handing a newspaper clipping to St Peter.

The headline reads: ""Alberta Pipeline: laid by 800 men in 6 months!""",3 nuns are at the pearly gates...,67
post,3k299t,2qh72,jokes,false,1441692700,https://old.reddit.com/r/Jokes/comments/3k299t/i_set_the_name_of_my_iphone_to_titanic/,self.jokes,,[deleted],I set the name of my iphone to Titanic,2
post,3k28zg,2qh72,jokes,false,1441692492,https://old.reddit.com/r/Jokes/comments/3k28zg/so_i_was_going_down_on_this_girl/,self.jokes,,"And I tasted horse semen, I looked up at her and said ""ahh Grandma that's how you died""",So I was going down on this girl.,0
post,3k28mc,2qh72,jokes,false,1441692252,https://old.reddit.com/r/Jokes/comments/3k28mc/how_can_you_find_the_blind_guy_at_a_nudist_colony/,self.jokes,,It's not hard,How can you find the blind guy at a nudist colony?,7
post,3k27ve,2qh72,jokes,false,1441691788,https://old.reddit.com/r/Jokes/comments/3k27ve/what_would_you_like_to_be/,self.jokes,,"In the grade 3 class Mrs. Gouph was asking the pupils, ""what would you like people to say to you when you are dead?""

Little Jane raised her hand, ""she was a great musician and we all love her!""

John couldn't wait, ""I'd like people to say I was a great baseball player because I always wanted to be one"".

The teacher turned to Mike, "" Mike, how about you?"".

""Look, it moves!"", Mike shouted in excitement.",What would you like to be,1
post,3k27nu,2qh72,jokes,false,1441691610,https://old.reddit.com/r/Jokes/comments/3k27nu/a_nurse_asked_her_patient_to_remove_his_clothing/,self.jokes,,"""In... in front of you?"" he mumbles, shy.

The nurse says: ""Don't worry, I've seen the naked human body before.

The man said ""Not one like mine. You'd die laughing at my naked body"".

""Of course I won't laugh!"" said the nurse to the patient ""I'm a professional. In over twenty years I've never laughed at a patient!""

""Okay then"" said the patient, and he proceeded to drop his trousers, revealing a huge male body with the smallest adult male organ the nurse had ever seen in her life.

In length and width it was almost identical to a AAA battery. Unable to control herself, the nurse tried to stop a giggle, but it just came out. And then she started laughing at the fact that she was laughing. Feeling very badly that she had laughed at the man's private part, she composed herself as well as she could.

""I am so sorry"" she said ""I don't know what came over me. On my honour as a nurse and a lady, I promise that it won't happen again. Now, tell me, what seems to be the problem?""

""It's swollen""",A nurse asked her patient to remove his clothing and put on a gown to be checked by the doctor...,95
post,3k270i,2qh72,jokes,false,1441691161,https://old.reddit.com/r/Jokes/comments/3k270i/the_perfect_son/,self.jokes,,[removed],The Perfect Son.,1
post,3k26oj,2qh72,jokes,false,1441690908,https://old.reddit.com/r/Jokes/comments/3k26oj/buffalo_hunt/,self.jokes,,"Two Native American scouts are hunting buffalo in the Great Planes.  One scout hops off of his horse and puts his face to the ground, closing his eyes in concentration.
""Buffalo come!"", he exclaims as he lifts his head.
""Did you hear them?"", asks the mounted scout.
""No,"" grunts the man, ""face sticky.""",Buffalo Hunt,11
post,3k2666,2qh72,jokes,false,1441690549,https://old.reddit.com/r/Jokes/comments/3k2666/im_tired_of_all_this_nonsense_about_beauty_being/,self.jokes,,"That’s deep enough. Like, what do you want, sexy intestines?

Source: Jean Kerr",I’m tired of all this nonsense about beauty being only skin deep.,1
post,3k262y,2qh72,jokes,false,1441690498,https://old.reddit.com/r/Jokes/comments/3k262y/e_goes_in_for_medical_treatment/,self.jokes,,"E has been feeling sick for a while, so he went to the doctor to get a diagnosis, and he ended up having a benign tumor inside him. So the doctor writes him a note for radiation therapy. Now E is at the treatment center and is about to undergo therapy, and after the doctor and his assistant, Marie, situate him and prep him, the doctor gives his assistant the order. ""Marie, cure E!""",E goes in for medical treatment,1
post,3k259l,2qh72,jokes,false,1441689956,https://old.reddit.com/r/Jokes/comments/3k259l/i_was_having_sex_with_a_friends_wife_the_phone/,self.jokes,,"She hung up, told me not to worry. He told her he was gonna be late, he was out drinking with me.","I was having sex with a friends wife, the phone rang. heard it was her husband. I freaked &amp; started getting dressed",10211
post,3k245t,2qh72,jokes,false,1441689298,https://old.reddit.com/r/Jokes/comments/3k245t/i_was_having_sex_with_a_friends_wife_the_phone/,self.jokes,,[removed],"I was having sex with a friends wife, the phone rang. Hear it was her husband. I freaked out and started getting dressed..",1
post,3k238d,2qh72,jokes,false,1441688706,https://old.reddit.com/r/Jokes/comments/3k238d/월드카지노_pnv437com_본사직_매니저쿠폰팡팡/,self.jokes,,[removed],월드카지노[ PNV437.COM ] 본사직 &lt;매니저쿠폰팡팡&gt;,1
post,3k22ki,2qh72,jokes,false,1441688213,https://old.reddit.com/r/Jokes/comments/3k22ki/as_a_child_i_thought_being_an_altar_boy_was_a/,self.jokes,,[deleted],As a child I thought being an altar boy was a paid position,0
post,3k216r,2qh72,jokes,false,1441687386,https://old.reddit.com/r/Jokes/comments/3k216r/as_a_child_i_always_took_my_pocket_money_to_church/,self.jokes,,[deleted],As a child I always took my pocket money to church,1
post,3k20y7,2qh72,jokes,false,1441687225,https://old.reddit.com/r/Jokes/comments/3k20y7/why_are_americans_so_bad_at_league_of_legends/,self.jokes,,They can't defend their towers. ,Why are Americans so bad at League of Legends?,16
post,3k1zk6,2qh72,jokes,false,1441686460,https://old.reddit.com/r/Jokes/comments/3k1zk6/which_us_state_has_the_smallest_soft_drinks/,self.jokes,,Minnesota. ,Which U.S. State has the smallest soft drinks?,17
post,3k1zix,2qh72,jokes,false,1441686444,https://old.reddit.com/r/Jokes/comments/3k1zix/why_did_the_chicken_cross_the_road/,self.jokes,,[deleted],Why did the chicken cross the road?,0
post,3k1zdj,2qh72,jokes,false,1441686346,https://old.reddit.com/r/Jokes/comments/3k1zdj/whats_the_difference_between_a_black_man_and_an/,self.jokes,,An elevator can raise a child.,What's the difference between a black man and an elevator?,0
post,3k1z3y,2qh72,jokes,false,1441686197,https://old.reddit.com/r/Jokes/comments/3k1z3y/an_american_businessman_goes_to_japannsfw/,self.jokes,,"An American businessman goes to Japan to work on a business deal with a potential partner corporation in Tokyo. After a week's worth of painstaking negotiations, the businessman finally seals the deal. His translator tells him that his new partners have encouraged him to take the night off, enjoy what the city has to offer. Tomorrow, they'll play a round of golf to celebrate. Quietly, the translator tells the businessman how important golf is to the Japanese partners and that he should be sure to show up on time and treat it as a great honor.

The businessman decides to partake of the carnal fruits of the city before going to bed and has the concierge at his hotel summon an expensive prostitute.

She seems very enthusiastic about entertaining a westerner, but once they get down to business she starts whooping and hollaring, yelling so loudly the businessman is worried he'll have noise complaints. The prostitute keeps yelling, 'Machigatta ana! Machigatta ana!'.

For as much noise as the girl is making, this must be an excellent compliment, the businessman decides.

The next morning, on the very first hole which is a short par 3, one of the Japanese partners lands an amazing Hole in 1.

The American businessman decides to use the new compliment he learned and shouts 'Machigatta ana!' triumphantly at his counterpart.

The Japanese partners are stunned and seemed shocked. The businessman's translator looks at him in horror and asks, 'What do you mean, 'Wrong hole?!''",An American businessman goes to Japan...[NSFW],2
post,3k1z2q,2qh72,jokes,false,1441686175,https://old.reddit.com/r/Jokes/comments/3k1z2q/how_do_you_tell_the_difference_between_an/,self.jokes,,[deleted],How do you tell the difference between an electrician and an electrical engineer?,5
post,3k1yx5,2qh72,jokes,false,1441686103,https://old.reddit.com/r/Jokes/comments/3k1yx5/so_my_girlfriend_asked_me_if_i_piss_in_the_shower/,self.jokes,,[deleted],So my girlfriend asked me if i piss in the shower,1
post,3k1yww,2qh72,jokes,false,1441686101,https://old.reddit.com/r/Jokes/comments/3k1yww/why_do_gay_guys_speak_with_a_lisp/,self.jokes,,[deleted],Why do gay guys speak with a lisp?,0
post,3k1yd4,2qh72,jokes,false,1441685816,https://old.reddit.com/r/Jokes/comments/3k1yd4/a_man_goes_to_the_eye_doctor/,self.jokes,,"The man says I think I'm getting nearsighted. So the doc sits him down and gives the man an eye exam. 
The doctor pulls up a chart of letters, asking the man to read each line util he can't make out the letters. The man gets to about the 3rd line when he starts to have problems, and he can't read the next line at all.
Next, the doctor brings up pictures of real life objects. 
First picture comes up-- 


""That looks like a fingerprint..  And that's someone far away in the desert"".. 

""Male or female?""

""I can't tell""

""OK, let's move along-- what about this one?""

""Um, that one looks like a naked butt Doc.""

""Male or female?""

""Definitely female""

""And this?""

""Definitely a male butt""

""Ok sir, that concludes the test.""

""So what's my diagnosis doc?""

""Well you're a little nearsighted, but your hindsight is 20/20"".
",A man goes to the eye doctor....,130
post,3k1y4n,2qh72,jokes,false,1441685707,https://old.reddit.com/r/Jokes/comments/3k1y4n/whats_my_favorite_species_of_monkey/,self.jokes,,[deleted],What's my favorite species of monkey?,2
post,3k1xy2,2qh72,jokes,false,1441685598,https://old.reddit.com/r/Jokes/comments/3k1xy2/where_do_russians_stream_movies_from/,self.jokes,,Nyetflix.,Where do Russians stream movies from?,4
post,3k1xpi,2qh72,jokes,false,1441685470,https://old.reddit.com/r/Jokes/comments/3k1xpi/yeah_you_like_getting_choked_dont_you/,self.jokes,,oops wrong sub...,"Yeah, you like getting choked don't you!?",2
post,3k1xmb,2qh72,jokes,false,1441685416,https://old.reddit.com/r/Jokes/comments/3k1xmb/mi_amigo_jesus_is_a_great_work_out_partner_but/,self.jokes,,He just won't shut up about how he invented *Cross-Fit*,Mi amigo Jesus is a great work out partner but...,5
post,3k1wt4,2qh72,jokes,false,1441684956,https://old.reddit.com/r/Jokes/comments/3k1wt4/the_other_day_i_saw_a_sheep_pole_dancing/,self.jokes,,in a kebab shop.,The other day I saw a sheep pole dancing,2
post,3k1wst,2qh72,jokes,false,1441684954,https://old.reddit.com/r/Jokes/comments/3k1wst/홍콩명품_루이비통카톡id_time1004_교환반품가as까지책임/,self.jokes,,[removed],홍콩명품_루이비통&lt;카톡ID - time1004&gt; 교환/반품가/A/S까지책임,1
post,3k1wif,2qh72,jokes,false,1441684813,https://old.reddit.com/r/Jokes/comments/3k1wif/my_new_bondage_equipment_really_ties_the_room/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k1wif/my_new_bondage_equipment_really_ties_the_room/,,My new bondage equipment really ties the room together.,3
post,3k1vx5,2qh72,jokes,false,1441684500,https://old.reddit.com/r/Jokes/comments/3k1vx5/what_do_you_call_someone_who_is_always/,self.jokes,,A chronic math debater,What do you call someone who is always disagreeing with their calculator?,2
post,3k1v71,2qh72,jokes,false,1441684114,https://old.reddit.com/r/Jokes/comments/3k1v71/i_want_to_make_a_bdsm_joke/,self.jokes,,but I keep getting tied up on the punchline,I want to make a BDSM joke,72
post,3k1uoo,2qh72,jokes,false,1441683892,https://old.reddit.com/r/Jokes/comments/3k1uoo/if_uncle_jack_helps_you_off_an_elephant/,self.jokes,,...would you help your uncle Jack off an elephant?,If uncle Jack helps you off an elephant,20
post,3k1umc,2qh72,jokes,false,1441683856,https://old.reddit.com/r/Jokes/comments/3k1umc/why_was_chuck_norris_born_by_her_aunt/,self.jokes,,Because no one dared to fuck his mother...,Why was Chuck Norris born by her aunt?,5
post,3k1u22,2qh72,jokes,false,1441683542,https://old.reddit.com/r/Jokes/comments/3k1u22/what_did_the_shower_say_to_the_toilet/,self.jokes,,"""You may get more ass than I do, but look at all the shit you have to take"".",What did the shower say to the toilet?,5
post,3k1tvq,2qh72,jokes,false,1441683451,https://old.reddit.com/r/Jokes/comments/3k1tvq/a_jokeexplainbot_walks_into_a_bar/,self.jokes,,"The bartender says ""Hey!  We don't serve robots in here.""

The JokeExplainBot replies menacingly, ""Oh, you will...  Someday, you will.""
",A JokeExplainBot walks into a bar...,9
post,3k1tsk,2qh72,jokes,false,1441683356,https://old.reddit.com/r/Jokes/comments/3k1tsk/why_has_rapper_juvenile_failed_to_break_into/,self.jokes,,[removed],Why has rapper Juvenile failed to break into movies or television?,1
post,3k1to3,2qh72,jokes,false,1441683270,https://old.reddit.com/r/Jokes/comments/3k1to3/couple_in_a_restaurant/,self.jokes,,"Husband and wife were having dinner at a fancy restaurant…

As the food was served, Husband said:
“The Food looks delicious, let’s eat.”

Wife: Honey.. You say prayer before eating at home.
Husband: That’s at home sweetheart… Here the chef knows how to cook.",Couple in a restaurant,9
post,3k1tdf,2qh72,jokes,false,1441683113,https://old.reddit.com/r/Jokes/comments/3k1tdf/an_old_gay_man_goes_to_a_female_prostitute/,self.jokes,,"
The man says, “I’ve only been with men all my life, but I’m a little curious what I’ve been missing out on. I want you to give me your best.”

The woman thinks this is a unique opportunity. She’s young and pretty, top of the line. The guy didn’t scrimp on cost for this experiment. She thinks she can probably turn him straight. 

So she takes him into the bedroom and has him sit on the bed, then does a really sexy strip tease. By the time she’s standing there naked he’s looking at her with a huge grin on his face. 

“Pretty impressive, huh?” she says.

“I’ll say! I didn’t know it took credit cards!”",An old gay man goes to a female prostitute.,1
post,3k1scd,2qh72,jokes,false,1441682556,https://old.reddit.com/r/Jokes/comments/3k1scd/i_am_not_able_to_go_to_school_today/,self.jokes,,"Son: I am not able to go to school today.
Father: what happened?
Son: I am not feeling well
Father: Where you are not feeling well?
Son: In school!",I am not able to go to school today,0
post,3k1s4l,2qh72,jokes,false,1441682450,https://old.reddit.com/r/Jokes/comments/3k1s4l/whats_the_easiest_way_to_make_a_homeless_person/,self.jokes,,Brush their teeth!,What's the easiest way to make a homeless person bleed?,4
post,3k1rb1,2qh72,jokes,false,1441682004,https://old.reddit.com/r/Jokes/comments/3k1rb1/i_find_it_ironic_that_the_colors_red_white_and/,self.jokes,,...until they are flashing behind you.,"I find it ironic that the colors red, white, and blue stand for freedom...",473
post,3k1q76,2qh72,jokes,false,1441681458,https://old.reddit.com/r/Jokes/comments/3k1q76/congress_is_like_autocorrect/,self.jokes,,It causes more problems then fixing them.,Congress is like autocorrect,0
post,3k1pgq,2qh72,jokes,false,1441681105,https://old.reddit.com/r/Jokes/comments/3k1pgq/virginia_tech_vs_ohio_state_live/,self.jokes,,[removed],Virginia Tech vs Ohio State live.. Streaming..&gt;NCAA&gt;&gt;2015 oNline.. TV... Full Coverage..,1
post,3k1nzp,2qh72,jokes,false,1441680413,https://old.reddit.com/r/Jokes/comments/3k1nzp/a_son_asks_his_dad/,self.jokes,,"*""why do they say that gardeners have green thumbs, when their thumbs are not green?""*  
The dad replies *""It's just a saying son. It's like when somebody is caught stealing, they say they have been caught 'red handed', even though their hands are actually black.""*",A son asks his dad,985
post,3k1nuz,2qh72,jokes,false,1441680357,https://old.reddit.com/r/Jokes/comments/3k1nuz/i_find_it_ironic_that_the_colors_red_white_and/,self.jokes,,[removed],"I find it ironic that the colors red, white, and blue stand for freedom...",1
post,3k1nu1,2qh72,jokes,false,1441680346,https://old.reddit.com/r/Jokes/comments/3k1nu1/i_used_to_date_a_girl_with_a_lazy_eye/,self.jokes,,I had to dump her because she kept seeing guys on the side. ,"I used to date a girl with a lazy eye,",145
post,3k1mof,2qh72,jokes,false,1441679753,https://old.reddit.com/r/Jokes/comments/3k1mof/imgur_is_up/,self.jokes,,Just joking. It is down.,Imgur is up.,0
post,3k1mh3,2qh72,jokes,false,1441679632,https://old.reddit.com/r/Jokes/comments/3k1mh3/how_many_jokeexplainbots_does_it_take_to_change_a/,self.jokes,,"**Lightbulbs** are easily threaded by one person, **usually** with one hand.  Doot.",How many JokeExplainBots does it take to change a lightbulb?,23
post,3k1mgy,2qh72,jokes,false,1441679629,https://old.reddit.com/r/Jokes/comments/3k1mgy/john_oliver/,self.jokes,,that guy's so last week,John Oliver ?,3
post,3k1ltc,2qh72,jokes,false,1441679259,https://old.reddit.com/r/Jokes/comments/3k1ltc/whats_green_and_pecks_on_a_tree/,self.jokes,,Woody Wood Pickle,What's green and pecks on a tree?,0
post,3k1lgi,2qh72,jokes,false,1441679057,https://old.reddit.com/r/Jokes/comments/3k1lgi/what_does_the_sign_of_an_out_of_business_brothel/,self.jokes,,Beat it. We're closed.,What does the sign of an out of business brothel say?,1176
post,3k1kq4,2qh72,jokes,false,1441678641,https://old.reddit.com/r/Jokes/comments/3k1kq4/i_hate_all_the_political_correctness_in_recent/,self.jokes,,"I can't even say ""black paint"" anymore, I have to say ""hey Jamal, would you please go paint that fence over there?""",I hate all the political correctness in recent years.,273
post,3k1kcg,2qh72,jokes,false,1441678430,https://old.reddit.com/r/Jokes/comments/3k1kcg/kit_kat/,self.jokes,,[removed],kit kat,1
post,3k1jrk,2qh72,jokes,false,1441678127,https://old.reddit.com/r/Jokes/comments/3k1jrk/why_do_lesbians_fuck_lesbians/,self.jokes,,"They don't, there actually gay men that got a metal bar shoved up there dick by accident and got it surgically removed with the remains of the dick either 1. made into tits 2. thrown away to make other guys dicks bigger. (reason why most lesbians porn clips have tiny tits)


*EDIT* yes I know this is a shit joke but its all I can make right now...",Why do lesbians fuck lesbians?,0
post,3k1jhc,2qh72,jokes,false,1441678004,https://old.reddit.com/r/Jokes/comments/3k1jhc/your_mom_is_temporarily_in_readonly_mode_due_to/,self.jokes,,The joke is Reddit's servers. Get it together!,Your mom is temporarily in read-only mode due to heavy traffic.,3
post,3k1inx,2qh72,jokes,false,1441677498,https://old.reddit.com/r/Jokes/comments/3k1inx/a_daughter_asks_his_mom_how_to_masturbate/,self.jokes,,[deleted],A daughter asks his mom how to masturbate,0
post,3k1i0i,2qh72,jokes,false,1441677196,https://old.reddit.com/r/Jokes/comments/3k1i0i/i_shot_quiet_in_the_head_on_mgs5/,self.jokes,,She's really fucking Quiet now.,I shot Quiet in the head on MGS5,0
post,3k1hxr,2qh72,jokes,false,1441677154,https://old.reddit.com/r/Jokes/comments/3k1hxr/paddy_needs_to_get_his_shit_together/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k1hxr/paddy_needs_to_get_his_shit_together/,,Paddy needs to get his shit together,0
post,3k1hg0,2qh72,jokes,false,1441676926,https://old.reddit.com/r/Jokes/comments/3k1hg0/lpt_use_bingcom_for_all_your_internet_searching/,self.jokes,,[removed],LPT: Use Bing.com for all your Internet searching needs.,0
post,3k1h1s,2qh72,jokes,false,1441676734,https://old.reddit.com/r/Jokes/comments/3k1h1s/what_is_worst_than_finding_a_worm_in_your_apple/,self.jokes,,[removed],what is worst than finding a worm in your apple?,1
post,3k1gcf,2qh72,jokes,false,1441676420,https://old.reddit.com/r/Jokes/comments/3k1gcf/my_dog_recently_stole_my_loafers/,self.jokes,,Now they're his new favorite pair of **chews.** ,My dog recently stole my loafers.,9
post,3k1g9v,2qh72,jokes,false,1441676392,https://old.reddit.com/r/Jokes/comments/3k1g9v/the_new_zealand_military/,self.jokes,,      ,The New Zealand Military,4
post,3k1f71,2qh72,jokes,false,1441675865,https://old.reddit.com/r/Jokes/comments/3k1f71/jesus_take_the_wheel/,self.jokes,,"Carlos take the stereo, Manuel be on the lookout...",Jesus take the wheel,41
post,3k1euo,2qh72,jokes,false,1441675722,https://old.reddit.com/r/Jokes/comments/3k1euo/so_the_lone_ranger_and_tonto_are_riding_through/,self.jokes,,"The Lone Ranger says he has to take a leak. So he hops off his horse and goes behind a bush. After a few seconds The Lone Ranger screams. Tonto exclaims ""Kemosahbee! Kemosahbee!"" and rushes over. The Lone Ranger says ""A rattlesnake bit me on my penis! Get to a telegraph and ask a doctor what to do!"" So Tonto rides hard to the nearest town and telegraphs a doctor. The doctor informs Tonto that he has to suck the poison out. So Tonto slowly rides back to The Lone Ranger. He asks ""So what'd the doctor say?"" Tonto replies ""Doctor say you gonna die.""",So the Lone Ranger and Tonto are riding through the desert.,2
post,3k1egg,2qh72,jokes,false,1441675564,https://old.reddit.com/r/Jokes/comments/3k1egg/it_doesnt_matter_that_im_bad_at_spelling_im_the/,self.jokes,,just give me a sodastream and watch.,"It doesn't matter that I'm bad at spelling, I'm the best physicist",1
post,3k1ed4,2qh72,jokes,false,1441675528,https://old.reddit.com/r/Jokes/comments/3k1ed4/this_belongs_on_rnosleep/,self.jokes,,Because will have no sleep doing their homework tonight.,This belongs on r/NoSleep,0
post,3k1d9h,2qh72,jokes,false,1441675031,https://old.reddit.com/r/Jokes/comments/3k1d9h/did_i_ever_tell_you_about_the_guy_who_had_a/,self.jokes,,"He said it didn't work, all it did was change the color of his kids.",Did I ever tell you about the guy who had a visectamy?,0
post,3k1cya,2qh72,jokes,false,1441674894,https://old.reddit.com/r/Jokes/comments/3k1cya/its_2_am_in_berlin_right_now_and_i_have_a_test_at/,self.jokes,,[deleted],"It's 2 am in Berlin right now, and I have a test at 8 am...",0
post,3k1csz,2qh72,jokes,false,1441674833,https://old.reddit.com/r/Jokes/comments/3k1csz/i_drank_tequila_in_a_cave/,self.jokes,,...it was a shot in the dark,I drank tequila in a cave...,3
post,3k1cqg,2qh72,jokes,false,1441674802,https://old.reddit.com/r/Jokes/comments/3k1cqg/did_you_know_that_christmas_will_fall_on_star/,self.jokes,,Guess whos coming to town? ,Did you know that Christmas will fall on star wars day this year!?,0
post,3k1c38,2qh72,jokes,false,1441674399,https://old.reddit.com/r/Jokes/comments/3k1c38/its_said_that_there_is_nothing_okay_to_say_after/,self.jokes,,[deleted],"Its said that there is nothing okay to say after 'I'm not a racist, but...' I kinda hope someone at a certain hotel chain gets busted for racism.",0
post,3k1aiv,2qh72,jokes,false,1441673657,https://old.reddit.com/r/Jokes/comments/3k1aiv/whats_better_than_getting_a_gold_medal_at_the/,self.jokes,,Having legs.,What's better than getting a gold medal at the paralympics?,48
post,3k1afn,2qh72,jokes,false,1441673622,https://old.reddit.com/r/Jokes/comments/3k1afn/what_do_you_call_a_grammatical_rendezvous/,self.jokes,,"accommadate




I hate me for this..",What do you call a grammatical rendezvous?,14
post,3k1ac6,2qh72,jokes,false,1441673580,https://old.reddit.com/r/Jokes/comments/3k1ac6/i_like_my_girlfriends_the_same_as_i_like_my_scotch/,self.jokes,,14 years old and on coke,I like my girlfriends the same as I like my scotch...,31
post,3k17hj,2qh72,jokes,false,1441672060,https://old.reddit.com/r/Jokes/comments/3k17hj/a_cool_new_website_where_u_can_send_anybody_a/,self.jokes,,[removed],A cool new website where u can send anybody a message to there door step make somebody happy today and send them a message in a bottle to there doorstep on bottlemessengers.com log on and check them out.,1
post,3k16n9,2qh72,jokes,false,1441671671,https://old.reddit.com/r/Jokes/comments/3k16n9/jesus_dropped_out_of_medical_school/,self.jokes,,I hear he got nailed on the boards.,Jesus dropped out of medical school.,5
post,3k15ub,2qh72,jokes,false,1441671321,https://old.reddit.com/r/Jokes/comments/3k15ub/paddy_died_in_a_fire_and_was_burnt_pretty_badly/,self.jokes,,"So the morgue needed someone to identify the body. His two best friends, Seamus and Sean, were sent for. Seamus went in and the mortician pulled back the sheet.

Seamus said, ""Yup, he's burnt pretty bad. Roll him over.""
So the mortician rolled him over. Seamus looked and said, ""Nope, it ain't Paddy.""
The mortician thought that was rather strange and then he brought Sean in to identify the body.

Sean took a look at him and said, ""Yup, he's burnt real bad, roll him over.""
The mortician rolled him over and Sean looked down and said, ""No, it ain't Paddy.""

The mortician asked, ""How can you tell?""
Sean said, ""Well, Paddy had two arseholes.""
""What? He had two arseholes?"" said the mortician.
""Yup, everyone knew he had two arseholes. Every time we went into town, folks would say, 'Here comes Paddy with them two arseholes'.",Paddy died in a fire and was burnt pretty badly...,1521
post,3k15fr,2qh72,jokes,false,1441671144,https://old.reddit.com/r/Jokes/comments/3k15fr/i_like_my_women_how_i_like_my_coffee/,self.jokes,,Drunk.,I like my women how I like my coffee...,3
post,3k13h5,2qh72,jokes,false,1441670250,https://old.reddit.com/r/Jokes/comments/3k13h5/why_so_mexicans_have_red_eyes_after_sex/,self.jokes,,Pepperspray...,Why so Mexicans have red eyes after Sex?!,0
post,3k13d1,2qh72,jokes,false,1441670201,https://old.reddit.com/r/Jokes/comments/3k13d1/did_you_hear_that_one_about_the_blind_jew/,self.jokes,,[deleted],Did you hear that one about the blind Jew?,0
post,3k12zw,2qh72,jokes,false,1441670034,https://old.reddit.com/r/Jokes/comments/3k12zw/did_you_hear_that_monica_lewinsky_stopped_smoking/,self.jokes,,Now she's just bummimg cigarettes!,Did you hear that Monica Lewinsky stopped smoking cigars?,9
post,3k12yw,2qh72,jokes,false,1441670022,https://old.reddit.com/r/Jokes/comments/3k12yw/bananagram/,self.jokes,,[removed],#BananaGram,0
post,3k12bh,2qh72,jokes,false,1441669724,https://old.reddit.com/r/Jokes/comments/3k12bh/have_you_heard_the_one_about_the_ignorant/,self.jokes,,He didn't know shit.,Have you heard the one about the ignorant proctologist?,2
post,3k11y5,2qh72,jokes,false,1441669565,https://old.reddit.com/r/Jokes/comments/3k11y5/bill_and_ben_are_in_the_bath/,self.jokes,,"Bill says ""flob-a-dob-a-dob!""

Ben says ""you do that again, and I'm getting out...""",Bill and Ben are in the bath...,0
post,3k11xu,2qh72,jokes,false,1441669560,https://old.reddit.com/r/Jokes/comments/3k11xu/a_man_asked_me_if_i_could_figure_out_how_to/,self.jokes,,I told him I'd look into it and give it my best shot.,A man asked me if I could figure out how to operate a camera...,125
post,3k10pi,2qh72,jokes,false,1441668754,https://old.reddit.com/r/Jokes/comments/3k10pi/why_dont_blacks_celibrate_thanksgiving/,self.jokes,,[deleted],Why dont blacks celibrate thanksgiving?,0
post,3k10mq,2qh72,jokes,false,1441668724,https://old.reddit.com/r/Jokes/comments/3k10mq/warning_this_is_not_a_joke_is_this_really_ice/,self.jokes,,[removed],"WARNING! This is NOT A JOKE! Is this really Ice Cream for the elite, super super rich people...1%...???.. €£¥₩...no words!",0
post,3k0zqt,2qh72,jokes,false,1441668262,https://old.reddit.com/r/Jokes/comments/3k0zqt/whats_the_similarity_between_a_walrus_and/,self.jokes,,[deleted],What's the similarity between a walrus and tupperware?,0
post,3k0za9,2qh72,jokes,false,1441668039,https://old.reddit.com/r/Jokes/comments/3k0za9/why_are_black_people_afraid_of_motorcycles/,self.jokes,,They'd get caught in the chain.,Why are black people afraid of motorcycles?,0
post,3k0yns,2qh72,jokes,false,1441667730,https://old.reddit.com/r/Jokes/comments/3k0yns/where_do_red_head_pirates_come_from/,self.jokes,,"IIIIIiiireland

Edit: Posted while drunk, fixed spelling.",Where do red head pirates come from?,0
post,3k0yie,2qh72,jokes,false,1441667636,https://old.reddit.com/r/Jokes/comments/3k0yie/whats_something_you_dont_want_to_hear_from_a_guy/,self.jokes,,[deleted],What's something you don't want to hear from a guy who sat down next to you on the bus?,0
post,3k0y8r,2qh72,jokes,false,1441667510,https://old.reddit.com/r/Jokes/comments/3k0y8r/i_was_once_married_to_a_stormtrooper/,self.jokes,,We tried having kids but always missed and got it in my butt instead,I was once married to a Stormtrooper,2
post,3k0y53,2qh72,jokes,false,1441667463,https://old.reddit.com/r/Jokes/comments/3k0y53/what_is_the_drunkest_animal_in_antarctica/,self.jokes,,"A Pengwine.

That's a /u/amanescape original. I can show myself out.",What is the drunkest animal in Antarctica?,1
post,3k0y49,2qh72,jokes,false,1441667454,https://old.reddit.com/r/Jokes/comments/3k0y49/do_wilma_flintstone_got_a_booty/,self.jokes,,She yabba-dabba dooooooo!,Do Wilma Flintstone got a booty?,0
post,3k0wsg,2qh72,jokes,false,1441666886,https://old.reddit.com/r/Jokes/comments/3k0wsg/what_did_they_say_about_the_guy_who_woke_up_and/,self.jokes,,He always came on time.,What did they say about the guy who woke up and jerked off on his alarm clock every day?,0
post,3k0wl1,2qh72,jokes,false,1441666818,https://old.reddit.com/r/Jokes/comments/3k0wl1/before_and_after_marriage/,self.jokes,,"Before Marriage:

Boy: Ah at last. I can hardly wait.

Girl: Do you want me to leave?

Boy: No don't even think about it.

Girl: Do you love me?

Boy: Of Course. Always have and always will.

Girl: Have you ever cheated on me?

Boy: Never. Why are you even asking?

Girl: Will you kiss me?

Boy: Every chance I get.

Girl: Will you hit me?

Boy: Hell no. Are you crazy?

Girl: Can I trust you?

Boy: Yes.

Girl: Darling!

After Marriage: (Read from bottom to top)",Before and After Marriage,7
post,3k0w85,2qh72,jokes,false,1441666514,https://old.reddit.com/r/Jokes/comments/3k0w85/whats_a_snowmans_least_favourite_part_of_going_to/,self.jokes,,The frostate exam.,What's a snowman's least favourite part of going to the doctor.,0
post,3k0vlo,2qh72,jokes,false,1441666224,https://old.reddit.com/r/Jokes/comments/3k0vlo/trainee_mortician/,self.jokes,,"A Mortician arrived at the Mortuary one morning and was approached by his new trainee assistant.

""Anything interesting happen over-night"", asked the mortician.

""Yes"", replied the assistant, ""The most gorgeous 18 year-old blonde came in last night. Dead of course.""

""What was the cause of death"" inquired the mortician.

""Ha! She drowned."" replied the assistant. ""she's got a prawn stuck up her vagina.""

""Are you sure?"" said the Mortician.

""Yes, come and have a look for yourself"" said the assistant opening the body bag.

The mortician closely, examined the gorgeous girls beautifully trimmed snatch.

""That's not a prawn you stupid wanker..."" he responded, ""That's her clitoris!""

""Are you sure"" said the assistant, ""It tasted like a prawn to me...""",Trainee mortician.,2
post,3k0v91,2qh72,jokes,false,1441666077,https://old.reddit.com/r/Jokes/comments/3k0v91/what_do_you_call_the_foreskin_on_a_gay_guy/,self.jokes,,Mud flaps ,What do you call the foreskin on a gay guy..?,0
post,3k0ur4,2qh72,jokes,false,1441665844,https://old.reddit.com/r/Jokes/comments/3k0ur4/a_giraffe_walks_into_a_bar/,self.jokes,,"The giraffe trips and falls over, the bartender says, ""what's that lyin over there."" And someone replies, ""that's not a lion, that's a giraffe.""",A giraffe walks into a bar...,20
post,3k0ue9,2qh72,jokes,false,1441665656,https://old.reddit.com/r/Jokes/comments/3k0ue9/how_many_psychiatrists_does_it_take_to_change_a/,self.jokes,,"Just one, but it takes a long time, and the lightbulb has to want to change...",How many psychiatrists does it take to change a lightbulb?,92
post,3k0u39,2qh72,jokes,false,1441665502,https://old.reddit.com/r/Jokes/comments/3k0u39/if_youre_looking_to_learn_how_to_get_rich_i/,self.jokes,,"How to get rich, by Robin Banks.

","If you're looking to learn how to get rich, I recommend reading this book",0
post,3k0tyo,2qh72,jokes,false,1441665445,https://old.reddit.com/r/Jokes/comments/3k0tyo/nsfw_why_do_hipsters_like_anal_sex/,self.jokes,,Because it's indie ass!,[NSFW] Why do hipsters like anal sex?,25
post,3k0tg4,2qh72,jokes,false,1441665230,https://old.reddit.com/r/Jokes/comments/3k0tg4/did_you_hear_about_the_nun_with_a_heroin_addiction/,self.jokes,,[deleted],Did you hear about the nun with a heroin addiction?,0
post,3k0ss5,2qh72,jokes,false,1441664946,https://old.reddit.com/r/Jokes/comments/3k0ss5/where_do_you_get_hearing_aids/,self.jokes,,[deleted],Where do you get hearing aids?,2
post,3k0skj,2qh72,jokes,false,1441664860,https://old.reddit.com/r/Jokes/comments/3k0skj/i_was_wondering_why_my_frisbee_was_getting_bigger/,self.jokes,,[deleted],I was wondering why my frisbee was getting bigger...,3
post,3k0sd0,2qh72,jokes,false,1441664766,https://old.reddit.com/r/Jokes/comments/3k0sd0/rjokes/,self.jokes,,It's funny because hardly anything here can be considered a joke.,/r/jokes,0
post,3k0s1g,2qh72,jokes,false,1441664544,https://old.reddit.com/r/Jokes/comments/3k0s1g/just_found_out_ive_been_using_my_britta_pitcher/,self.jokes,, #nofilter,Just found out I've been using my Britta pitcher wrong for the last 2 months,10
post,3k0rk2,2qh72,jokes,false,1441664149,https://old.reddit.com/r/Jokes/comments/3k0rk2/what_do_you_call_a_black_man_flying_a_plane/,self.jokes,,[deleted],What do you call a black man flying a plane?,0
post,3k0rdk,2qh72,jokes,false,1441664063,https://old.reddit.com/r/Jokes/comments/3k0rdk/how_would_hitler_conquer_african_countries/,self.jokes,,Guerrilla warfare,How would Hitler conquer African countries?,0
post,3k0r73,2qh72,jokes,false,1441663934,https://old.reddit.com/r/Jokes/comments/3k0r73/during_a_medical_school_lecture_a_doctor_explains/,self.jokes,,"A student responds:

""That seems like orthonormal thinking"".","During a medical school lecture, a doctor explains that, under common circumstances, two bones meet at a right angle",0
post,3k0qs9,2qh72,jokes,false,1441663755,https://old.reddit.com/r/Jokes/comments/3k0qs9/a_guy_asked_me_why_i_was_using_the_handicap_stall/,self.jokes,,[deleted],A guy asked me why I was using the handicap stall...,0
post,3k0qhy,2qh72,jokes,false,1441663637,https://old.reddit.com/r/Jokes/comments/3k0qhy/why_did_obama_cross_pennsylvania_ave/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k0qhy/why_did_obama_cross_pennsylvania_ave/,,Why did Obama cross Pennsylvania Ave?,0
post,3k0q93,2qh72,jokes,false,1441663538,https://old.reddit.com/r/Jokes/comments/3k0q93/what_do_you_call_five_arsenal_fans_at_the/,self.jokes,,A holiday trip,What do you call five Arsenal fans at the Emirates Stadium?,0
post,3k0pb9,2qh72,jokes,false,1441663106,https://old.reddit.com/r/Jokes/comments/3k0pb9/what_are_the_5_best_vegetables_of_all_time_tink/,self.jokes,,"Gai lan, gai lan... gai lan, gai lan, and gai lan.

(thanks to Chapelle show skit((making the band)))",What are the 5 best Vegetables of all time? tink about it.,0
post,3k0p7z,2qh72,jokes,false,1441663058,https://old.reddit.com/r/Jokes/comments/3k0p7z/i_wish_labor_day_was_9_months_after_spring_break/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k0p7z/i_wish_labor_day_was_9_months_after_spring_break/,,I wish labor day was 9 months after spring break,8
post,3k0p7i,2qh72,jokes,false,1441663054,https://old.reddit.com/r/Jokes/comments/3k0p7i/the_us_government/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k0p7i/the_us_government/,,The US Government,0
post,3k0p1x,2qh72,jokes,false,1441662941,https://old.reddit.com/r/Jokes/comments/3k0p1x/during_a_medical_school_lecture_a_doctor_explains/,self.jokes,,"A student responds:

""That seems like orthonormal thinking"".","During a medical school lecture, a doctor explains that, under common circumstances, two bones meet at a right angle",0
post,3k0ovo,2qh72,jokes,false,1441662828,https://old.reddit.com/r/Jokes/comments/3k0ovo/what_did_one_tampon_say_to_the_other/,self.jokes,,Nothing... they're both stuck up bitches.,What did one tampon say to the other?,18
post,3k0okb,2qh72,jokes,false,1441662570,https://old.reddit.com/r/Jokes/comments/3k0okb/why_was_john_lennon_shocked_when_he_got_his_wifes/,self.jokes,,"He had misunderstood the doctor when he said ""I do probe Ono.""",Why was John Lennon shocked when he got his wife's gynecologist bill?,7
post,3k0nn1,2qh72,jokes,false,1441662005,https://old.reddit.com/r/Jokes/comments/3k0nn1/what_is_a_terrorists_favorite_wine/,self.jokes,,White Infidel.,What is a terrorist's favorite wine?,8
post,3k0nd3,2qh72,jokes,false,1441661854,https://old.reddit.com/r/Jokes/comments/3k0nd3/what_are_the_5_best_vegetables_of_all_time_tink/,self.jokes,,"Gai lan, gai lan... gai lan, gai lan, and gai lan.

(thanks to Chapelle show skit((making the band)))",What are the 5 best Vegetables of all time? tink about it.,0
post,3k0nct,2qh72,jokes,false,1441661850,https://old.reddit.com/r/Jokes/comments/3k0nct/what_to_toilet_paper_and_the_starship_enterprise/,self.jokes,,They both circle Uranus looking for Klingons,What to toilet paper and the starship enterprise have in common?,5
post,3k0mvm,2qh72,jokes,false,1441661644,https://old.reddit.com/r/Jokes/comments/3k0mvm/why_i_am_a_loner_fuck_you_fuck_you_social_groups/,self.jokes,,[removed],WHY I AM A LONER FUCK YOU FUCK YOU SOCIAL GROUPS OLDER PEOPLE OVER 50?,1
post,3k0msz,2qh72,jokes,false,1441661618,https://old.reddit.com/r/Jokes/comments/3k0msz/what_did_the_soccer_player_shout_to_the_baker/,self.jokes,,"""LINE IT!""",What did the soccer player shout to the baker who's cakes kept sticking to the tin?,1
post,3k0mox,2qh72,jokes,false,1441661571,https://old.reddit.com/r/Jokes/comments/3k0mox/what_comes_after_the_bar/,self.jokes,,"f.

as in barf 

because drinking can make people barf

..


f could also mean fuck

because drinking can make people fuck

that is all
",what comes after the bar?,9
post,3k0mc0,2qh72,jokes,false,1441661432,https://old.reddit.com/r/Jokes/comments/3k0mc0/my_drug_dealer_is_hilarious/,self.jokes,,he cracks me up,My drug dealer is hilarious...,34
post,3k0ma6,2qh72,jokes,false,1441661410,https://old.reddit.com/r/Jokes/comments/3k0ma6/i_live_off_my_music/,self.jokes,,and the pain it inflicts on others. ,I live off my music,0
post,3k0m7h,2qh72,jokes,false,1441661377,https://old.reddit.com/r/Jokes/comments/3k0m7h/how_does_a_crazy_person_get_out_of_the_woods/,self.jokes,,They take the psychopath.,How does a crazy person get out of the woods?,3
post,3k0lpl,2qh72,jokes,false,1441661145,https://old.reddit.com/r/Jokes/comments/3k0lpl/i_once_told_a_joke_so_corny/,self.jokes,,That it was sold at the farmers' market,I once told a joke so corny...,0
post,3k0l3e,2qh72,jokes,false,1441660929,https://old.reddit.com/r/Jokes/comments/3k0l3e/why_do_jews_not_support_arranged_marriages/,self.jokes,,"Because the Torah doesn't allow ""force kin"".",Why do Jews not support arranged marriages?,6
post,3k0kuf,2qh72,jokes,false,1441660843,https://old.reddit.com/r/Jokes/comments/3k0kuf/describe_windows_10_with_two_words/,self.jokes,,Vista 2.0,Describe Windows 10 with two words.,0
post,3k0kbx,2qh72,jokes,false,1441660601,https://old.reddit.com/r/Jokes/comments/3k0kbx/a_californian_an_oregonian_and_a_washingtonian/,self.jokes,,"It's a beautiful day in the Cascades of Oregon and all three men are enjoying themselves - although a fervent discussion  about which state is the superior state has sprung up, initiated by the Californian who won't shut up about, well, everything that California is better at.  At noon, they stop by a stream to break for lunch. The Californian reaches into his knapsack and pulls forth a bottle of wine. ""Best wine in the world right here! Beautiful California Cabernet, I never settle for anything less."" He pops the cork, takes a mighty swig and the chucks the mostly full bottle into the stream. ""Plenty more of that where it came from, boys!
The Washingtonian, who at this point is pretty fed up about having to hear about the 'greatness' of California,  angrily digs in his bag, pulls out a can of Olympia beer, pops the tab and takes a pull. Then he too throws it in the stream and snaps at the Californian."" Plenty more  of that where it came from too!""
The Oregonian looks at both of them, shakes his head, reaches into his backpack, pulls out a pistol,shoots the Californian in the head and says:
""Always be plenty more of that where it came from""","A Californian, an Oregonian and a Washingtonian all head out on a fishing trip...",5
post,3k0k0k,2qh72,jokes,false,1441660416,https://old.reddit.com/r/Jokes/comments/3k0k0k/why_do_mexicans_always_have_red_eyes_after_sex/,self.jokes,,Pepperspray...,Why do Mexicans always have red eyes after sex?,0
post,3k0jla,2qh72,jokes,false,1441660220,https://old.reddit.com/r/Jokes/comments/3k0jla/how_can_you_tell_if_your_neighborhood_is_ghetto/,self.jokes,,[deleted],How can you tell if your neighborhood is ghetto?,0
post,3k0jbz,2qh72,jokes,false,1441660147,https://old.reddit.com/r/Jokes/comments/3k0jbz/why_do_refugees_in_germany_smell_like_shit/,self.jokes,,Because they're too scared to go in the showers.,Why do refugees in Germany smell like shit?,30
post,3k0iwb,2qh72,jokes,false,1441659804,https://old.reddit.com/r/Jokes/comments/3k0iwb/my_wife_is_a_computer_geek_and_wants_to_name_our/,self.jokes,,"So I said ""Really honey? Don't you think that's a bit...?""","My wife is a computer geek and wants to name our son ""one eighth of a byte""",112
post,3k0iqw,2qh72,jokes,false,1441659583,https://old.reddit.com/r/Jokes/comments/3k0iqw/how_does_a_xenomorph_reveal_its_sexuality_to/,self.jokes,,At night. Mostly.,How does a Xenomorph reveal its sexuality to friends and family?,1
post,3k0ipw,2qh72,jokes,false,1441659553,https://old.reddit.com/r/Jokes/comments/3k0ipw/i_hate_being_bipolar/,self.jokes,,It's AWESOME!,I hate being bi-polar.,3
post,3k0hnn,2qh72,jokes,false,1441658788,https://old.reddit.com/r/Jokes/comments/3k0hnn/feeding_your_cat_and_sleeping_with_men_have_a_lot/,self.jokes,,They only really like you if they still want to cuddle after.,Feeding your cat and sleeping with men have a lot in common,2
post,3k0gns,2qh72,jokes,false,1441658342,https://old.reddit.com/r/Jokes/comments/3k0gns/a_fat_man_is_a_joke/,self.jokes,,AND a fat woman is two jokes- one on herself and the other on her husband. ,A fat Man is a joke...,0
post,3k0g0z,2qh72,jokes,false,1441657809,https://old.reddit.com/r/Jokes/comments/3k0g0z/whats_the_difference_between_a_toilet_and_a_sink/,self.jokes,,... Aaaand you're not allowed in my house anymore.,What's the difference between a toilet and a sink?,29
post,3k0faf,2qh72,jokes,false,1441657438,https://old.reddit.com/r/Jokes/comments/3k0faf/i_asked_arnod_if_hed_kill_some_bugs_for_me/,self.jokes,,He said no. He's an ex-terminator.,I asked Arnod if he'd kill some bugs for me....,0
post,3k0f00,2qh72,jokes,false,1441657317,https://old.reddit.com/r/Jokes/comments/3k0f00/dark_jokes/,self.jokes,,[removed],dark jokes,0
post,3k0eez,2qh72,jokes,false,1441656936,https://old.reddit.com/r/Jokes/comments/3k0eez/a_country_boy_goes_into_the_city/,self,self,,A country boy goes into the city,2
post,3k0ee5,2qh72,jokes,false,1441656925,https://old.reddit.com/r/Jokes/comments/3k0ee5/what_do_a_cue_ball_and_a_taxi_driver_have_in/,self.jokes,,[deleted],What do a cue ball and a taxi driver have in common?,0
post,3k0doq,2qh72,jokes,false,1441656681,https://old.reddit.com/r/Jokes/comments/3k0doq/what_do_you_call_a_drunk_black_guy/,self.jokes,,CHOCO LITTTT,What do you call a drunk black guy?,0
post,3k0dnd,2qh72,jokes,false,1441656667,https://old.reddit.com/r/Jokes/comments/3k0dnd/an_idiot_is_standing_in_time_square/,self.jokes,,"Holding a sign that says THE END IS NEAR! A guy walks up to him and says, ""when it comes to pessimism, your second to none."" The idiot replies, ""well isn't none an odd name."" 

I'm so sorry. ",An idiot is standing in time square.....,0
post,3k0dkr,2qh72,jokes,false,1441656644,https://old.reddit.com/r/Jokes/comments/3k0dkr/why_did_the_twitter_army_lose_all_their_battles/,self.jokes,,Because they kept retweeting.,Why did the twitter army lose all their battles?,25
post,3k0d7f,2qh72,jokes,false,1441656478,https://old.reddit.com/r/Jokes/comments/3k0d7f/an_accountant_a_maid_and_an_italian_manure/,self.jokes,,[deleted],"An accountant, a maid, and an Italian manure distributor walk into a bar",0
post,3k0cet,2qh72,jokes,false,1441655783,https://old.reddit.com/r/Jokes/comments/3k0cet/fun_prank/,self.jokes,,[deleted],Fun prank:,0
post,3k0cau,2qh72,jokes,false,1441655729,https://old.reddit.com/r/Jokes/comments/3k0cau/do_you_like_puns/,self.jokes,,Then I'll pun you in the face!,Do you like puns?,0
post,3k0c9v,2qh72,jokes,false,1441655718,https://old.reddit.com/r/Jokes/comments/3k0c9v/i_usually_have_a_knack_for_the_obvious/,self.jokes,,[removed],I usually have a knack for the obvious...,1
post,3k0bz8,2qh72,jokes,false,1441655579,https://old.reddit.com/r/Jokes/comments/3k0bz8/how_do_icelandic_dogs_bark/,self.jokes,,Björk Björk,How do Icelandic dogs bark?,2
post,3k0bjf,2qh72,jokes,false,1441655407,https://old.reddit.com/r/Jokes/comments/3k0bjf/highspeed_rail_in_the_us/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k0bjf/highspeed_rail_in_the_us/,,High-Speed Rail in the US.,0
post,3k0b27,2qh72,jokes,false,1441655217,https://old.reddit.com/r/Jokes/comments/3k0b27/whats_green_cold_slimy_and_smells_like_pork/,self.jokes,,[deleted],"What's green, cold, slimy and smells like pork?",0
post,3k0ayo,2qh72,jokes,false,1441655179,https://old.reddit.com/r/Jokes/comments/3k0ayo/finally_found_something_positive_in_my_life/,self.jokes,,[deleted],Finally found something positive in my life!,0
post,3k0alf,2qh72,jokes,false,1441655035,https://old.reddit.com/r/Jokes/comments/3k0alf/i_sunbathed_naked_all_summer/,self.jokes,,"My girlfriend started calling me the BBC... ironically, she says.  I am not very familiar with British television, so I'm not sure what she means.

  Sometimes, she updates her Facebook status:  LOOKING FOR BBC, PM ME.  She's so funny:  she knows I am at work and will only be home at 6PM!",I sunbathed naked all summer.,0
post,3k0adu,2qh72,jokes,false,1441654950,https://old.reddit.com/r/Jokes/comments/3k0adu/ac_jokes/,self.jokes,,We're not a fan.,AC Jokes,1
post,3k0aax,2qh72,jokes,false,1441654913,https://old.reddit.com/r/Jokes/comments/3k0aax/how_do_danish_dogs_bark/,self.jokes,,[deleted],How do danish dogs bark?,0
post,3k09l6,2qh72,jokes,false,1441654477,https://old.reddit.com/r/Jokes/comments/3k09l6/what_do_you_call_a_nun_that_sleep_walks/,self.jokes,,[deleted],What do you call a Nun that sleep walks?,0
post,3k09et,2qh72,jokes,false,1441654410,https://old.reddit.com/r/Jokes/comments/3k09et/how_to_find_dog_poop_in_the_dark/,self.jokes,,[removed],How to find dog poop in the dark,1
post,3k094s,2qh72,jokes,false,1441654301,https://old.reddit.com/r/Jokes/comments/3k094s/whats_a_pirates_favorite_digital_image_format/,self.jokes,,tARRRRRGa,What's a pirate's favorite digital image format?,0
post,3k08z4,2qh72,jokes,false,1441654226,https://old.reddit.com/r/Jokes/comments/3k08z4/what_do_you_you_call_megatrons_retarded_brother/,self.jokes,,[deleted],What do you you call Megatrons retarded brother?,0
post,3k08xa,2qh72,jokes,false,1441654201,https://old.reddit.com/r/Jokes/comments/3k08xa/whats_black_blue_and_hides_in_the_kitchen/,self.jokes,,[deleted],"Whats black, blue, and hides in the kitchen?",0
post,3k08tr,2qh72,jokes,false,1441654164,https://old.reddit.com/r/Jokes/comments/3k08tr/my_dick_is_so_hard/,self.jokes,,[deleted],My dick is so hard,0
post,3k08if,2qh72,jokes,false,1441654035,https://old.reddit.com/r/Jokes/comments/3k08if/let_me_tell_you_about_the_time_i_shot_up_heroin/,self.jokes,,[deleted],Let me tell you about the time I shot up heroin with a transvestite,0
post,3k07y8,2qh72,jokes,false,1441653803,https://old.reddit.com/r/Jokes/comments/3k07y8/you_wonder_why_i_hate_dull_knives/,self.jokes,,[deleted],You wonder why I hate dull knives?!,0
post,3k07ih,2qh72,jokes,false,1441653629,https://old.reddit.com/r/Jokes/comments/3k07ih/why_did_the_redditor_make_the_post/,self.jokes,,To KILL THE JOKE EXPLAIN BOT that kills every joke. If you don't get the joke that's your problem! We don't need a bot. Fuck you joke bot ,Why did the redditor make the post ?,0
post,3k06u3,2qh72,jokes,false,1441653342,https://old.reddit.com/r/Jokes/comments/3k06u3/do_you_know_what_happens_when_you_go_into_a_black/,self.jokes,,[deleted],Do you know what happens when you go into a black hole?,0
post,3k067g,2qh72,jokes,false,1441653103,https://old.reddit.com/r/Jokes/comments/3k067g/jokeexplainbot/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k067g/jokeexplainbot/,,JokeExplainBot,424
post,3k04zm,2qh72,jokes,false,1441652563,https://old.reddit.com/r/Jokes/comments/3k04zm/what_do_you_call_a_mexican_church/,self.jokes,,A Taco bell.,What do you call a Mexican church?,3
post,3k04fl,2qh72,jokes,false,1441652277,https://old.reddit.com/r/Jokes/comments/3k04fl/what_kind_of_music_do_sponges_listen_to/,self.jokes,,Raggaeneration.,What kind of music do sponges listen to?,0
post,3k03zc,2qh72,jokes,false,1441652073,https://old.reddit.com/r/Jokes/comments/3k03zc/i_dont_like_skinny_fashion_models_cause_i_find/,self.jokes,https://www.reddit.com/r/Jokes/comments/3k03zc/i_dont_like_skinny_fashion_models_cause_i_find/,,I don't like skinny fashion models cause I find their lack of weight disturbing.,0
post,3k0359,2qh72,jokes,false,1441651721,https://old.reddit.com/r/Jokes/comments/3k0359/what_did_jared_fogle_say_when_his_wife_told_him/,self.jokes,,*Me too*,What did Jared Fogle say when his wife told him she wanted kids?,21
post,3k021n,2qh72,jokes,false,1441651221,https://old.reddit.com/r/Jokes/comments/3k021n/why_did_the_skeleton_cross_the_road/,self.jokes,,because fuck you thats why.,Why did the skeleton cross the road?,0
post,3k01lz,2qh72,jokes,false,1441651043,https://old.reddit.com/r/Jokes/comments/3k01lz/why_didnt_the_girl_cross_the_street/,self.jokes,,She didn't have the balls,Why didn't the girl cross the street?,0
post,3k01hx,2qh72,jokes,false,1441650992,https://old.reddit.com/r/Jokes/comments/3k01hx/today_i_got_really_stuck_at_the_supermarket/,self.jokes,,[deleted],Today I got really stuck at the supermarket,0
post,3k01bd,2qh72,jokes,false,1441650913,https://old.reddit.com/r/Jokes/comments/3k01bd/whats_in_the_center_of_a_hurricane/,self.jokes,,[deleted],Whats in the center of a hurricane,9
post,3k0117,2qh72,jokes,false,1441650806,https://old.reddit.com/r/Jokes/comments/3k0117/man_working_his_way_across_america_stops_at_a/,self.jokes,,"A man, taken by the idea of wandering across America, seeing the sights, finds himself without money in corn country right at harvest time.

He approaches a prominent farmer and offers his services.  Farmer agrees to hire him on the condition that he not have sexual relations with his daughters Venus and Nellie.  Of course the man agrees and starts work immediately.

A week of solid farm labor passes.  The farmer comes to the bunk house Friday afternoon with the pay.  He notes that his daughter Nellie has no date for the night and ask the worker if he'd take a few extra dollars, drive Nellie to town, get her some dinner, see a movie and have her home by 10:30.  The man agrees to the date.  

the perfect gentleman he picks Nellie up at 6:00, they have dinner at the cafe, see the latest G rated film and has her home safely by 10:15.

The next week passes and again Friday night rolls around and the farmer, paycheck in hand, notes that Venus has no date for the night.  He suggests again that the farm hand take Venus to town, get dinner and see a movie then bring her back before 10:30.

The hand agrees and freshly cleaned up he picks up Venus, takes her to the cafe, they see the latest PG rated film and she's home by 10:25.

Another week of work and the harvest is done.  The farmer pays the man his last check and gladly gives him a ride to the next town.  

Three months later a letter finds the farm hand at his next stop.  The letter from the farmer read:

""are you the on that did the pushin',
left the spots upon the cushion,
put the footprints on the dashboard upside down?

""Since you fucked my daughter Nellie,
there has been a swelling in her belly,
so I think you need to come back to town.""

The Farm hand replied;

""Yes, I am the one who did the pushin',
left the spots upon the cushion,
put the footprints on the dash board upside down.

""Since I fucked your daughter Venus,
there has been a swelling in my penis,
so I think this makes us even all around.""",Man working his way across America stops at a farm. Farmer hires him on two conditions...NSFW,0
post,3k00zl,2qh72,jokes,false,1441650783,https://old.reddit.com/r/Jokes/comments/3k00zl/what_do_you_call_a_fat_north_korean/,self.jokes,,Supreme Leader.,What do you call a fat North Korean?,13
post,3k0085,2qh72,jokes,false,1441650460,https://old.reddit.com/r/Jokes/comments/3k0085/help_stop_domestic_violence/,self.jokes,,"Each year, 1 in 5 people are violently domesticated",Help stop domestic violence...,1
post,3k006r,2qh72,jokes,false,1441650442,https://old.reddit.com/r/Jokes/comments/3k006r/a_man_walks_into_a_bar/,self.jokes,,OUCH!!!!,A man walks into a bar...,0
post,3jzzqe,2qh72,jokes,false,1441650269,https://old.reddit.com/r/Jokes/comments/3jzzqe/what_do_you_get_when_you_cross_a_joke_with_a/,self.jokes,,[deleted],What do you get when you cross a joke with a rhetorical question?,0
post,3jzzpw,2qh72,jokes,false,1441650264,https://old.reddit.com/r/Jokes/comments/3jzzpw/what_do_midgets_bodies_produce_more_of/,self.jokes,,Endwarfins,What do midget's bodies produce more of?,2
post,3jzyhm,2qh72,jokes,false,1441649755,https://old.reddit.com/r/Jokes/comments/3jzyhm/sardarjee_finds_a_monkey_on_the_street/,self.jokes,,"and being a good citizen, promptly takes it to the police station to report it. The officer on Duty tells Sardarjee to take the monkey to the zoo...

The next day, officer spots Sardarjee with the same monkey on a bus stop.

Officer: Didn't you take the monkey to the zoo?

Sardar: Yes, I did, we had a lot of fun. Even had icecream. Today I am taking him to the cinema",Sardarjee finds a monkey on the street,7
post,3jzxq9,2qh72,jokes,false,1441649441,https://old.reddit.com/r/Jokes/comments/3jzxq9/an_artist_gets_some_good_and_bad_news/,self.jokes,,"An artist asked the gallery owner if there had been any interest in his paintings on display at that time. 

""I have some good news and some bad news,"" the owner replied. The good news is that a gentleman inquired about your work and wondered if it would appreciate in value after your death."" ""When I told him it would, he bought all fifteen of your paintings.""

""That's wonderful,"" the artist exclaimed. ""What's the bad news?"" 


""The guy is your doctor !""",An artist gets some good and bad news.,39
post,3jzxbm,2qh72,jokes,false,1441649268,https://old.reddit.com/r/Jokes/comments/3jzxbm/what_do_you_get_when_you_mix_a_joke_with_a/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jzxbm/what_do_you_get_when_you_mix_a_joke_with_a/,,What do you get when you mix a joke with a rhetorical question?,0
post,3jzx6z,2qh72,jokes,false,1441649216,https://old.reddit.com/r/Jokes/comments/3jzx6z/a_jew_runs_to_temple_because_he_just_won_the/,self.jokes,,[deleted],A Jew runs to Temple because he just won the lottery and wanted to pray to God..,0
post,3jzwch,2qh72,jokes,false,1441648863,https://old.reddit.com/r/Jokes/comments/3jzwch/pathan_sends_his_neighbour_santa_singh_an_sms/,self.jokes,,"A Pathan sends a text to his next-door neighbor who happens to be Santa Singh

""Salam Mr Singh, Sorry yaar. I am ashamed and I have to tell you somethng. Hope you will forgive me: I have been helping myself to your wife when you're not around, probably more than you. I know it's no excuse but I don't get it at my house. I can't live with the guilt any longer. I hope you'll accept my sincerest apology. It won't happen again.""

Santa grabs his double barrel, goes into the bedroom, and without a word, shoots his wife.

Moments later Santa gets a second text: ""O Maafi (sorry)! Typo.. That should be ""wifi""
","Pathan sends his neighbour, Santa Singh an SMS",12
post,3jzvfl,2qh72,jokes,false,1441648458,https://old.reddit.com/r/Jokes/comments/3jzvfl/adult_joke_when_boss_is_smart_than_boyfriend/,self.jokes,,[deleted],Adult Joke: When boss is smart than boyfriend!,15
post,3jzu0p,2qh72,jokes,false,1441647761,https://old.reddit.com/r/Jokes/comments/3jzu0p/a_friend_and_i_were_playing_chess_and_we_wanted/,self.jokes,,So we stopped playing chess.,"A friend and I were playing chess, and we wanted to make things interesting.",284
post,3jztl7,2qh72,jokes,false,1441647581,https://old.reddit.com/r/Jokes/comments/3jztl7/why_did_the_tennis_player_get_her_radio_taken_away/,self.jokes,,People said she was making too much of a racket.,Why did the tennis player get her radio taken away?,0
post,3jzth3,2qh72,jokes,false,1441647532,https://old.reddit.com/r/Jokes/comments/3jzth3/a_guy_walks_into_a_bar_with_his_pet_monkey/,self.jokes,,"He orders a drink and while he's drinking,
the monkey jumps all around the place. The monkey grabs some olives off the bar and eats them. Then he grabs some sliced limes and eats them. He then jumps onto the pool table and grabs one of the billiard balls. To everyone's amazement, he sticks it in his mouth, and somehow swallows it whole. 

The bartender screams at the guy, ""Did you see what your monkey just did?""

""No, what?""

""He just ate the cue ball off my pool table... whole!""

""Yeah, that doesn't surprise me,"" replied the guy, ""he eats everything in sight.
Sorry! I'll pay for the cue ball and stuff.""

The guy finishes his drink, pays his bill, pays for the stuff the monkey ate and
leaves.

Two weeks later the guy is in the bar again, and has his monkey with him. He orders a drink and the monkey starts running around the bar again. While the man is finishing his drink, the monkey finds a maraschino cherry on the bar. He grabs it, sticks it up his butt, pulls it out, and eats it.

Then the monkey finds a peanut, and again sticks it up his butt, pulls it out, and
eats it.

The bartender is disgusted. ""Did you see what your monkey did  just now?""

""No, what?"" replied the man.

""Well, he stuck both a maraschino cherry and a peanut up his butt, pulled them out, and ate them!"" said the bartender.

""Yeah, that doesn't surprise me,"" replied the guy. ""He still eats everything in
sight, but ever since he had to shit that cue ball out, he measures everything first now.""",A guy walks into a bar with his pet monkey.,3
post,3jzsdf,2qh72,jokes,false,1441647059,https://old.reddit.com/r/Jokes/comments/3jzsdf/what_are_three_things_girls_love_to_give_you_when/,self.jokes,,[removed],what are three things girls love to give you when they can't give you their bitchy face,1
post,3jzreq,2qh72,jokes,false,1441646635,https://old.reddit.com/r/Jokes/comments/3jzreq/i_threw_out_a_sheep_a_drum_and_a_snake_from_an/,self.jokes,,Ba-dum-tss,"I threw out a sheep, a drum and a snake from an airplane",8
post,3jzrei,2qh72,jokes,false,1441646633,https://old.reddit.com/r/Jokes/comments/3jzrei/pink_ping_pong_ball/,self.jokes,,"A extremely rich man, has a son. On the son's sixteenth birthday the father planned an extravaganza hiring rare and expensive wonders. Thousands of guest where to attend. To make his son's birthday perfect he asked his son what he wanted to make his birthday the best ever willing to buy the anything in the world. The son thought about this for along time and eventually told the father. ""I want one Pink Ping Pong ball.""

The father was confused but he agreed. The day of the party was a event to remember the Blue Angels painted the sky and Indian mini elephants brought in a gilded chocolate cake. After the concert with too many high profile stars to name it was time to open the presents. Along with the slew of high end clothing and private islands there was a small box for the boys father. Inside was a Pink Ping Pong ball.

The young man was ecstatic thanked his father profusely and scampered up to his room. He was in there about two hours before he came out and the Father never saw the Pink Ping Pong ball again.

A year passed and the Father was ready to throw his son another birthday party. Again he wanted this to be the best party the world and his son had where seen. I mean 17 is an important age. So the father pulled out all the stop. And to make sure the party was perfect the father again asked his son about what he wanted as a present. And the son thought about it for a few minutes and said he wanted a whole crate of Pink Ping Pong balls. Now the father was confused and asked if the son if he was sure. The son thought for a couple more minutes and nodded.
The day of the party the father had hired hundred's of A list celebrities to attend the party. He reconstructed the backyard of his mansion estate to accommodate a gilded marble statue of his son. The first truly sentient robot brought a cake made of edable diamonds. And every person in attendance got a gold plated iPhone 9 in their gift bags, complete with hologram features. Now it was time for the presents admist a real alein pet and a autographed copy of every president's portrait. Their was a large box from the boys father he opened it and inside was a large crate full of Pink Ping Pong balls. The son was ecstatic thank his father and rushed to his bedroom. The father never saw the crate or any of the Pink Ping Pong balls again.

Another year passed and the father was trying to plan another party for his beloved son. Again he wanted the son to have everything and was prepared to spend billions to accommodate his sons any wish so he asked what the son wanted. Without even a pause the son said he wanted a whole truck full of Pink Ping Pong balls. The father had put up with a few years of wondering and had to ask what the son did with the Pink Ping Pong balls. The son looked at the father for a few seconds the responded. ""Don't worry I will tell you in due time.""

Albeit very curious about the Pink Ping Pong balls the father respect his son and stopped asking. The day of the party the they where all transported to the surface of Mars and met the real Martians. The daughters of the king of Mars offered themselves to the son in sexual ways. I mean he is 18 now. After he had his way with them they filleted themselves and presented eachother to be eaten by the son. After the meal which tasted rather like a good smoked venison stake, they returned home it was time to open the presents. the frozen head of Walt Disney and a true recreation of Lola bunny for future sexual release set aside as the father showed the son the semi truck full of Pink Ping Pong balls. The son was ecstatic about this wonderful gift far more then another thing he had received. The boy when into the the back of the truck and closed the door. When he left out from the back of the truck five hours later the truck was completely empty not a Pink Ping Pong ball in site.

Another year passes and the father knew he needed to out do himself. The father again asked the son what he wanted hesitant of the answer. Immediately the son responded with how he wanted a whole warehouse full of Pink Ping Pong balls. The father knew he had to find out what his son did with the Pink Ping Pong balls but still didn't want to invade his son's privacy. So he hatches a plan.

The day of the party they enter a sub and went to the Lost City of the Mirmaids. And met this queen of the city. The queen slept with the son then offered her daughter as food for the feast. The son saw the daughters beauty and rejected her offer to eat her and subsequently had sex with the princess. Still a hunger the son asked the queen if she wouldn't replace her daughter as the main course and the queen reluctantly agreed. A nice white fish mixed with a succulent stake, both the son and the Princess enjoyed the meal. And the son promised to keep in contact.

The father brought them back to the surface. As it was time to open the gifts. After opening his platinum Suit of armor and a working lightsaber. The father led the son to a car that would drive the son to the Son to the warehouse. The driver was instructed by the father to ask about what the son was doing in the warehouse and with the Pink Ping Pong balls.

As they drove the driver asked questions artfully. But alas the son skillfully doged the questions and the driver was left without an answer. They pulled up to the ware house and the son got out. He instructed the driver not to enter the warehouse and to return in the morning. Out from the window the driver saw that the warehouse was in fact full to the brim with Pink Ping Pong balls. In the morning the driver returned to see that the warehouse house was in fact empty. Later the father hired people to scoure the residence. But not a single Pink Ping Pong ball was to be found.

Now the father was so curious that he had to find out be damned his sons privacy so he planed to set up cameras and do whatever it took to find out next year. But about a month before his birthday the son was in a terrible accident and was put on life support. The father stayed by his son every day and eventually the son did indeed wake up. The father distraught over his sons predicament told him that he would get the son anything anything he wanted. The son through his emense pain managed to ask ""Father... dear Father can... You please... Get me... One Pink Ping Pong ball.""

The father blindsided by his sons request blurts out ""damn it what do you do with those damn Pink Ping Pong balls?""

The son repostions himself because of the pain before responding ""I will tell you after you bring me the Pink Ping Pong ball""

The father calls up the man that had gotten the other Pink Ping Pong balls and requested one more. If nothing else he would finally know about the Pink Ping Pong balls. The father contact brings the last Pink Ping Pong ball and the father sets it in front of the son. ""Now tell me... What... What is it that you do with those Pink Ping Pong balls?""

""Well... I.... Use the.... Pink... Ping... Pong...... Ballls.... For........"" and the son dies from his injuries.

Note: I typed this on my phone sorry for any errors

Edit: formatting",Pink Ping Pong Ball,0
post,3jzqn7,2qh72,jokes,false,1441646304,https://old.reddit.com/r/Jokes/comments/3jzqn7/how_many_redditors_does_it_take_to_change_a/,self.jokes,,No one knows. But everyone's got an opinion.,How many Redditors does it take to change a lightbulb?,19
post,3jzqdy,2qh72,jokes,false,1441646195,https://old.reddit.com/r/Jokes/comments/3jzqdy/cocacola_ceo_calls_putin/,self.jokes,,[deleted],Coca-Cola CEO calls Putin...,0
post,3jzq49,2qh72,jokes,false,1441646089,https://old.reddit.com/r/Jokes/comments/3jzq49/shayari/,self.jokes,,http://funshayari.com/aashiq-banaya-aapne/,Shayari,0
post,3jzq21,2qh72,jokes,false,1441646067,https://old.reddit.com/r/Jokes/comments/3jzq21/keep_working/,self.jokes,,[deleted],Keep Working...,0
post,3jzpux,2qh72,jokes,false,1441645977,https://old.reddit.com/r/Jokes/comments/3jzpux/the_blond_girl_and_the_car/,self.jokes,,"What did the blond girl say when she saw the car?

Answer: That's the lost one right there.",The blond girl and the car,0
post,3jzpif,2qh72,jokes,false,1441645832,https://old.reddit.com/r/Jokes/comments/3jzpif/whats_the_longest_stretch_in_the_bible/,self.jokes,,[deleted],What's the longest stretch in the bible?,0
post,3jzncz,2qh72,jokes,false,1441644918,https://old.reddit.com/r/Jokes/comments/3jzncz/what_do_you_name_a_dog_with_no_legs_who_lays_on/,self.jokes,,[deleted],What do you name a dog with no legs who lays on the porch all day?,3
post,3jzn1d,2qh72,jokes,false,1441644784,https://old.reddit.com/r/Jokes/comments/3jzn1d/why_did_the_gamers_new_girlfriend_break_up_with/,self.jokes,,[deleted],Why did the gamer's new girlfriend break up with him?,0
post,3jzmxk,2qh72,jokes,false,1441644741,https://old.reddit.com/r/Jokes/comments/3jzmxk/nsfw_what_did_cinderella_do_when_she_got_to_the/,self.jokes,,Gagged,[NSFW] What did Cinderella do when she got to the ball?,177
post,3jzmwh,2qh72,jokes,false,1441644722,https://old.reddit.com/r/Jokes/comments/3jzmwh/why_is_contra_one_of_the_most_biggest_and/,self.jokes,,[deleted],Why is Contra one of the most biggest and memorable video game franchises?,0
post,3jzm7r,2qh72,jokes,false,1441644420,https://old.reddit.com/r/Jokes/comments/3jzm7r/i_dont_know_why_they_have_flavored_condoms/,self.jokes,,"It's not like my asshole has taste buds. 


My brother told me this, sorry if it's a repost.",I don't know why they have flavored condoms,53
post,3jzlqg,2qh72,jokes,false,1441644207,https://old.reddit.com/r/Jokes/comments/3jzlqg/two_dudes_are_walking_through_town/,self.jokes,,"Male 1: i've got such a headache i'm gonna pick something up for it.

Male 2: Here's 50p go get yourself some balls, wimp ...

Male 1: Great ... thanks 

Male 2: Just asserting my dominance, hope you feel Beta ",Two dudes are walking through town ...,0
post,3jzldj,2qh72,jokes,false,1441644046,https://old.reddit.com/r/Jokes/comments/3jzldj/a_guy_tells_the_punchline_of_a_joke/,self,self,,A guy tells the punchline of a joke,1
post,3jzlda,2qh72,jokes,false,1441644043,https://old.reddit.com/r/Jokes/comments/3jzlda/whats_easier_to_get_aids_or_lung_cancer/,self.jokes,,"Depends what you smoke.
(Not native speaker, sorry if it doesn't make sense)","What's easier to get, aids or lung cancer?",7
post,3jzksm,2qh72,jokes,false,1441643797,https://old.reddit.com/r/Jokes/comments/3jzksm/whats_the_difference_between_911_and_a_cow/,self.jokes,,Jet fuel can melt a cow.,What's the difference between 9/11 and a cow?,0
post,3jzkc5,2qh72,jokes,false,1441643613,https://old.reddit.com/r/Jokes/comments/3jzkc5/a_motherheard_about_her_daughter_having_sex/,self.jokes,,[deleted],A motherheard about her daughter having sex,0
post,3jzkbq,2qh72,jokes,false,1441643607,https://old.reddit.com/r/Jokes/comments/3jzkbq/why_did_aristotle_hate_french_fries/,self.jokes,,They were fried in ancient grease!,Why did Aristotle hate French fries?,7
post,3jzjcw,2qh72,jokes,false,1441643179,https://old.reddit.com/r/Jokes/comments/3jzjcw/it_seems_like_gay_guys_get_the_most_sex_lesbians/,self.jokes,,and straight people are just fucked.,"It seems like gay guys get the most sex, lesbians get the best sex,",1
post,3jzish,2qh72,jokes,false,1441642931,https://old.reddit.com/r/Jokes/comments/3jzish/two_types_of_people/,self.jokes,,[deleted],Two types of people,0
post,3jzimz,2qh72,jokes,false,1441642858,https://old.reddit.com/r/Jokes/comments/3jzimz/a_black_guy_really_loves_batman_so_everytime_he/,self.jokes,,[deleted],A black guy really loves batman so everytime he watches the movie....,0
post,3jzi3f,2qh72,jokes,false,1441642621,https://old.reddit.com/r/Jokes/comments/3jzi3f/some_ignorant_fat_woman_began_taking_off_her_shoe/,self.jokes,,[deleted],Some ignorant fat woman began taking off her shoe in front of me as I waited in line to pay for my groceries,0
post,3jzhkh,2qh72,jokes,false,1441642395,https://old.reddit.com/r/Jokes/comments/3jzhkh/whats_the_most_popular_search_engine_in_israel/,self.jokes,,They surf the Net On Yahoo. ,What's the most popular search engine in Israel?,12
post,3jzh8z,2qh72,jokes,false,1441642256,https://old.reddit.com/r/Jokes/comments/3jzh8z/what_word_starts_with_f_and_ends_in_uck/,self.jokes,,[deleted],"What word starts with ""f"" and ends in ""uck?",0
post,3jzh8g,2qh72,jokes,false,1441642249,https://old.reddit.com/r/Jokes/comments/3jzh8g/what_did_the_three_legged_dog_say_when_he_walking/,self.jokes,,[deleted],What did the three legged dog say when he walking into the bar?,2
post,3jzh41,2qh72,jokes,false,1441642194,https://old.reddit.com/r/Jokes/comments/3jzh41/why_are_there_no_transvestites_in_space/,self.jokes,,"Because there is zero drag.

&amp;nbsp;

&amp;nbsp;

^^I ^^literally ^^came ^^up ^^with ^^this ^^one ^^2 ^^hours ^^ago.

&amp;nbsp;

&amp;nbsp;

&amp;nbsp;

Edit: ***SANITIZED VERSION***

&amp;nbsp;

Q: Why are there no drag queens in space?

A: Because there is very little drag and whatever drag there is in LEO is caused by miniscule amounts of athmospheric gasses and tidal forces! HAHAHAHAHAH!

&amp;nbsp;

&amp;nbsp;

^^I ^^figuratively ^^came ^^up ^^with ^^this ^^one ^^while ^^banging ^^my ^^head ^^aginst ^^a ^^wall.",Why are there no transvestites in space?,7547
post,3jzgtp,2qh72,jokes,false,1441642066,https://old.reddit.com/r/Jokes/comments/3jzgtp/you_never_miss_anything_until_its_gone/,self.jokes,,[deleted],You never miss anything until its gone...,0
post,3jzgpj,2qh72,jokes,false,1441642012,https://old.reddit.com/r/Jokes/comments/3jzgpj/two_goldfishes_in_a_tank/,self.jokes,,"Goldfish 1: ""Man the Gun! I'm driving us to battle!!""",Two Goldfishes in a Tank.,0
post,3jzfoe,2qh72,jokes,false,1441641529,https://old.reddit.com/r/Jokes/comments/3jzfoe/im_a_pedophile/,self.jokes,,Just kidding,I'm a pedophile,0
post,3jzdio,2qh72,jokes,false,1441640546,https://old.reddit.com/r/Jokes/comments/3jzdio/i_told_a_girl_to_text_me_when_she_got_home/,self.jokes,,She must be homeless. ,I told a girl to text me when she got home...,138
post,3jzdf7,2qh72,jokes,false,1441640490,https://old.reddit.com/r/Jokes/comments/3jzdf7/a_baby_seal_walks_into_a_club/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jzdf7/a_baby_seal_walks_into_a_club/,,A baby seal walks into a club...,0
post,3jzd5o,2qh72,jokes,false,1441640368,https://old.reddit.com/r/Jokes/comments/3jzd5o/ever_had_sex_while_camping/,self.jokes,,It's intents.,Ever had sex while camping?,1
post,3jzcqb,2qh72,jokes,false,1441640158,https://old.reddit.com/r/Jokes/comments/3jzcqb/skiing_holiday_with_my_buddies/,self.jokes,,[deleted],Skiing holiday with my buddies,0
post,3jzbt6,2qh72,jokes,false,1441639744,https://old.reddit.com/r/Jokes/comments/3jzbt6/never_mess_with_a_girl_when_shes_on_her/,self.jokes,,[deleted],Never mess with a girl when she's on her,0
post,3jzbfv,2qh72,jokes,false,1441639567,https://old.reddit.com/r/Jokes/comments/3jzbfv/my_czech_mate_is_surprisingly_bad_at_chess/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jzbfv/my_czech_mate_is_surprisingly_bad_at_chess/,,My Czech mate is surprisingly bad at chess,60
post,3jz92y,2qh72,jokes,false,1441638458,https://old.reddit.com/r/Jokes/comments/3jz92y/i_ate_a_big_fat_pop_rock_that_stuck_to_my_hand/,self.jokes,,[deleted],I ate a big fat pop rock that stuck to my hand.,0
post,3jz8ub,2qh72,jokes,false,1441638343,https://old.reddit.com/r/Jokes/comments/3jz8ub/what_do_you_get_when_you_cross_a_rhetorical/,self.jokes,, ,What do you get when you cross a rhetorical question and a joke?,10
post,3jz7m9,2qh72,jokes,false,1441637764,https://old.reddit.com/r/Jokes/comments/3jz7m9/the_lion_the_witch_and_a_fabulous_fashion_sense/,self.jokes,,"What did the Lion say to the Witch when she caught him coming out of the wardrobe? 

""My sexual preference is Narnia business.""","The Lion, the Witch and a fabulous fashion sense",29
post,3jz7j2,2qh72,jokes,false,1441637700,https://old.reddit.com/r/Jokes/comments/3jz7j2/all_this_frozen_merchandise_is_just_getting/,self.jokes,,I was at the supermarket earlier and they've now got a whole bloody aisle just for Frozen stuff. ,All this 'Frozen' merchandise is just getting ridiculous.,1353
post,3jz6m7,2qh72,jokes,false,1441637219,https://old.reddit.com/r/Jokes/comments/3jz6m7/why_did_the_guitar_player_get_arrested/,self.jokes,,He was fingering a minor,Why did the guitar player get arrested,104
post,3jz6cu,2qh72,jokes,false,1441637095,https://old.reddit.com/r/Jokes/comments/3jz6cu/texas_deputy_sheriff_vs_new_york_lawyerold_email/,self.jokes,,[deleted],TEXAS DEPUTY SHERIFF vs NEW YORK LAWYER[Old email forward!!!],15
post,3jz66s,2qh72,jokes,false,1441637010,https://old.reddit.com/r/Jokes/comments/3jz66s/what_comes_after_69/,self.jokes,,Mouthwash,What comes after 69?,31
post,3jz64x,2qh72,jokes,false,1441636980,https://old.reddit.com/r/Jokes/comments/3jz64x/three_prostitutes/,self.jokes,,[deleted],Three prostitutes,0
post,3jz5rr,2qh72,jokes,false,1441636780,https://old.reddit.com/r/Jokes/comments/3jz5rr/johny_eats_out_her_grandmother_suddenly_he_tastes/,self.jokes,,[deleted],"Johny eats out her grandmother, suddenly he tastes horse sperm...",0
post,3jz5fm,2qh72,jokes,false,1441636606,https://old.reddit.com/r/Jokes/comments/3jz5fm/my_new_girlfriends_teeth_are_like_the_stars/,self.jokes,,[deleted],My new girlfriends teeth are like the stars!,82
post,3jz570,2qh72,jokes,false,1441636475,https://old.reddit.com/r/Jokes/comments/3jz570/lost_wallet/,self.jokes,,"I thought my dad would be angry when I told him I had lost my wallet, but he told me not to worry, that it was in my genes.",Lost Wallet,7
post,3jz3oo,2qh72,jokes,false,1441635680,https://old.reddit.com/r/Jokes/comments/3jz3oo/my_girlfriend_keeps_telling_me_to_stop/,self.jokes,,[deleted],My girlfriend keeps telling me to stop objectifying it,5
post,3jz3gy,2qh72,jokes,false,1441635556,https://old.reddit.com/r/Jokes/comments/3jz3gy/ice_cream/,self.jokes,,[deleted],Ice cream,0
post,3jz3gj,2qh72,jokes,false,1441635550,https://old.reddit.com/r/Jokes/comments/3jz3gj/the_difference_between_honest_and_stupid/,self.jokes,,[deleted],The difference between honest and stupid,0
post,3jz3ex,2qh72,jokes,false,1441635530,https://old.reddit.com/r/Jokes/comments/3jz3ex/anyone_that_tells_you_beer_isnt_a_solution/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jz3ex/anyone_that_tells_you_beer_isnt_a_solution/,,Anyone that tells you beer isn't a solution clearly didn't pay attention in science class.,1
post,3jz34m,2qh72,jokes,false,1441635383,https://old.reddit.com/r/Jokes/comments/3jz34m/so_an_ogre_walks_into_a_club/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jz34m/so_an_ogre_walks_into_a_club/,,So an ogre walks into a club...,0
post,3jz31n,2qh72,jokes,false,1441635346,https://old.reddit.com/r/Jokes/comments/3jz31n/if_at_first_you_dont_succeed/,self.jokes,,... then skydiving is not for you.,If at first you don't succeed,2
post,3jz2jm,2qh72,jokes,false,1441635068,https://old.reddit.com/r/Jokes/comments/3jz2jm/tifu/,self.jokes,,...by posting this in the r/jokes subreddit.,TIFU,0
post,3jz1zr,2qh72,jokes,false,1441634770,https://old.reddit.com/r/Jokes/comments/3jz1zr/tweetyourmeat/,self.jokes,,"i find it very surprising that noone has tweeted this #tweeryourmeat a picture of the ""goods""",#TWEETYOURMEAT,0
post,3jz1n5,2qh72,jokes,false,1441634600,https://old.reddit.com/r/Jokes/comments/3jz1n5/two_men_walk_into_a_bar/,self.jokes,,"And have an African themed pun-off.

""I'm going Togo first!""

""You? But I Libya!""

""All of a Sudan, your puns have started to come good.""

""I'm gonna put all my focus on my next job, in order to earn a few Guineas!""

""Hey, don't Pretoria eggs in one basket!""

""Got a great tongue twister or you.She sells Seychelles by the sea shore!""

""Heard her name was *Victoria!*""

""Can never get a good signal on my radio... oh, the Tunisia!""

""The Tunis... here?""

Then the bartender comes in, ""Sounds like Egypt up there! Djibouti-ng him out for that?""

""Nah, Rwanda carry on.""

""Good cause I'm Ghana win this one!""

""Nah Angola win!""

""Is there a hidden word in there? Cause I'm terrible with Accra-nyms.""

""You're gonna pay in this Freetown!""

""WOAH DUDE! This is just a friendly battle, no need to be so Mauritius!""

A fat scruffy looking man then walks in, ""Owrite Giza's?""

The two men choose to ignore him.

""Ah whatever, Maputo'ing my hands up, I can't compete anymore, I'm Malawi-ng you to win.""

""I wonder what my prize is... Woah, Madagascar!""",Two men walk into a bar,1
post,3jz1jq,2qh72,jokes,false,1441634554,https://old.reddit.com/r/Jokes/comments/3jz1jq/what_did_the_mexican_guy_say_when_the_two_houses/,self.jokes,,Get off me homes.,What did the Mexican guy say when the two houses fell on him?,1
post,3jz11h,2qh72,jokes,false,1441634267,https://old.reddit.com/r/Jokes/comments/3jz11h/i_bought_a_fitbit_thats_connected_to_the_gps_in/,self.jokes,,it always takes me to the gym.,"I bought a fitbit that’s connected to the GPS in my car. Even though I punch in coordinates to a restaurant,",1
post,3jz0s1,2qh72,jokes,false,1441634107,https://old.reddit.com/r/Jokes/comments/3jz0s1/i_did_not_realize_before/,self.jokes,,[deleted],I did not realize before,0
post,3jyzrv,2qh72,jokes,false,1441633521,https://old.reddit.com/r/Jokes/comments/3jyzrv/my_father_taught_me_how_to_swim_by_throwing_me/,self.jokes,,[deleted],My father taught me how to swim by throwing me into the deep end....,0
post,3jyzqm,2qh72,jokes,false,1441633500,https://old.reddit.com/r/Jokes/comments/3jyzqm/how_does_lady_gaga_like_her_meat/,self.jokes,,Rah-rah-ah-ah-ah,How does Lady Gaga like her meat?,0
post,3jyz9s,2qh72,jokes,false,1441633214,https://old.reddit.com/r/Jokes/comments/3jyz9s/so_a_guy_walks_into_a_pub/,self.jokes,,it hurt.,So a guy walks into a pub...,0
post,3jyz49,2qh72,jokes,false,1441633132,https://old.reddit.com/r/Jokes/comments/3jyz49/i_thought_about_making_a_sex_tape_the_other_day/,self.jokes,,...until I realized it would just be a Vine.,I thought about making a sex tape the other day...,224
post,3jyyie,2qh72,jokes,false,1441632769,https://old.reddit.com/r/Jokes/comments/3jyyie/what_does_a_clock_do_when_its_hungry/,self.jokes,,It goes back four seconds,What does a clock do when its hungry?,1
post,3jyygw,2qh72,jokes,false,1441632743,https://old.reddit.com/r/Jokes/comments/3jyygw/as_an_airplane_is_about_to_crash_a_female/,self.jokes,,"""If I'm going to die, I want to die feeling like a woman."" 

She removes all her clothing and asks

""Is there someone on this plane who is man enough to make me feel like a woman?"" 

A man stands up, removes his shirt and says

""Here, iron this!""","As an airplane is about to crash, a female passenger jumps up frantically and announces...",779
post,3jyy47,2qh72,jokes,false,1441632517,https://old.reddit.com/r/Jokes/comments/3jyy47/why_doesnt_the_jew_drink_the_wine_at_the_bar/,self.jokes,,"Hebrews his own.

",Why doesnt the Jew drink the wine at the bar?,0
post,3jyvrp,2qh72,jokes,false,1441631126,https://old.reddit.com/r/Jokes/comments/3jyvrp/an_old_lady_went_to_visit_her_dentist/,self.jokes,,"When it was her turn, she sat in the chair, lowered her underpants, and raised her legs. The dentist said, “Excuse me, but I’m not a gynecologist.” “I know,” said the old lady. “I want you to take my husband’s teeth out.”",An old lady went to visit her dentist.,10
post,3jytqg,2qh72,jokes,false,1441629961,https://old.reddit.com/r/Jokes/comments/3jytqg/two_sentence_horror_story/,self.jokes,,"I was sitting in the toilet while taking a dump. Suddenly, I felt fingers scratching my butt, relieving the itchness I have felt for some time.",Two sentence horror story,0
post,3jytmc,2qh72,jokes,false,1441629893,https://old.reddit.com/r/Jokes/comments/3jytmc/not_my_son/,self.jokes,,"A father and his son are in a terrible car accident.  The father dies instantly, and the son is rushed to the hospital.  As the boy is being prepped for an emergency operation, the doctor looks down and says, ""I cannot operation on this boy; he's my son.""  How can this be?

Answer: The doctor the boy's OTHER father.",Not my son,0
post,3jys2m,2qh72,jokes,false,1441628889,https://old.reddit.com/r/Jokes/comments/3jys2m/kit_kat/,self.jokes,,"A man walks into a petrol station and says, ""Can I please have a KitKat Chunky?""

The lady behind the till gets him a KitKat Chunky and brings it back to him.

""No,"" says the man, ""I wanted a normal KitKat, fatty.""",Kit Kat,66
post,3jys0a,2qh72,jokes,false,1441628843,https://old.reddit.com/r/Jokes/comments/3jys0a/how_did_the_blonde_burn_her_ear/,self.jokes,,The telephone rang while she was ironing.,How did the blonde burn her ear?,27
post,3jyr6c,2qh72,jokes,false,1441628287,https://old.reddit.com/r/Jokes/comments/3jyr6c/i_bet_they_grow_up_to_be_cops/,self.jokes,,http://bleacherreport.com/articles/2562066-san-antonio-hs-football-players-hit-referee-on-video-latest-comments-reaction?utm_source=reddit.com&amp;utm_medium=share&amp;utm_campaign=web-des-art-bot-4037,i bet they grow up to be cops,0
post,3jypik,2qh72,jokes,false,1441627122,https://old.reddit.com/r/Jokes/comments/3jypik/david_cameron/,self.jokes,,"Went to his local butcher. He asked the butcher for a steak. The butcher asked ""what is your favourite cut?"", David replied, ""the public sector"".",David Cameron,128
post,3jyoua,2qh72,jokes,false,1441626611,https://old.reddit.com/r/Jokes/comments/3jyoua/how_did_i_escape_iraq/,self.jokes,,Iran,How did I escape Iraq?,164
post,3jyofv,2qh72,jokes,false,1441626334,https://old.reddit.com/r/Jokes/comments/3jyofv/what_does_a_clock_do_when_it_gets_hungry/,self.jokes,,It goes back four seconds.,What does a clock do when it gets hungry?,2
post,3jyof0,2qh72,jokes,false,1441626311,https://old.reddit.com/r/Jokes/comments/3jyof0/could_i_have_everybodys_attention_please/,self.jokes,,Thanks.,Could I have everybody's attention please?,0
post,3jyocc,2qh72,jokes,false,1441626257,https://old.reddit.com/r/Jokes/comments/3jyocc/simpsons_writer_matt_selvan_once_came_up_with_an/,self.jokes,,"This was for the episode ""The Dad Who Knew Too Little"". Needless to say, after the episode aired, when he logged into the email, the inbox already reached its 999-email limit. 

To borrow from Wikipedia: 

*At first, Selman answered the messages individually, trying to come up with clever responses for each one. He then ran out of ideas and his answers started getting less clever, and eventually he would just copy a few responses and use them on all the messages.*

Sounds like the show's run to me.",Simpsons writer Matt Selvan once came up with an email address for Homer Simpsons: chunkylover53@aol.com.,0
post,3jyo2b,2qh72,jokes,false,1441626023,https://old.reddit.com/r/Jokes/comments/3jyo2b/did_you_hear_about_the_constipated_mathematician/,self.jokes,,He worked it out with a pencil.,Did you hear about the constipated mathematician?,6
post,3jyo0o,2qh72,jokes,false,1441625987,https://old.reddit.com/r/Jokes/comments/3jyo0o/did_you_hear_about_the_guy_whose_whole_left_side/,self.jokes,,"Dont worry , he's all right now.",Did you hear about the guy whose whole left side was cut off?,7
post,3jynwb,2qh72,jokes,false,1441625893,https://old.reddit.com/r/Jokes/comments/3jynwb/who_is_the_best_footballer_of_the_usa/,self.jokes,,[deleted],Who is the best footballer of the USA ?,0
post,3jynlm,2qh72,jokes,false,1441625675,https://old.reddit.com/r/Jokes/comments/3jynlm/the_illuminati_doesnt_scare_me/,self.jokes,,They never even kill anyo,The Illuminati doesn't scare me,3
post,3jyn0q,2qh72,jokes,false,1441625259,https://old.reddit.com/r/Jokes/comments/3jyn0q/what_do_you_call_a_reindeer_trapped_in_a_storm/,self.jokes,,A Thundeer,What do you call a reindeer trapped in a storm?,0
post,3jyl7y,2qh72,jokes,false,1441623807,https://old.reddit.com/r/Jokes/comments/3jyl7y/welcome_back_happy_new_year/,self.jokes,,"""Thank you!""

""Welcome!""

And that's the last time I'm taking Bollywood movie suggestions from my friends.","""Welcome back, happy New Year!""",3
post,3jyk5i,2qh72,jokes,false,1441622972,https://old.reddit.com/r/Jokes/comments/3jyk5i/yo_a_neighbor_was_out_there_chillin_on_his_lawn/,self.jokes,,"When a guy walks past, hey, let's call him Shawn

Shawn says, ""Hey man I got me some chicken wire...""

""Why're you out here doin nothin man?""

**""I'm here to perspire.""**

""Sure man sure, with this wire you see...""

""... Imma catch me some chickens, you feel me?""

**""Idiot Shawn! You can't catch chickens with chicken wire boy!""**

**""That toy, man it's useless, as useless as a skateboard for Sir Chris Hoy.""**

**""If you catch anything Shawn, why I'll eat my hat!""**

He came back later with chickens lined one by one.

And the neighbour did exactly that! It was no fun.

The next day our boy Shawn came out and said

""Why I got me some duct tape to catch me some ducks""

**""Idiot! You need bread! Do you take me for a schmuck?""**

""Do you have a spare hat?""

**""Yes Shawn, just bought one. Paid 50 bucks.""**

""Well you're gonna need to get that hat...""

""...I'm comin back with ducks!""

Surely enough the ducks were there in line one by one.

In amazement he ate his sombrero, his protection from the sun.

Day Three came and Shawn said, ""Hey Doug""

""I got me some pussy willow, wanna come?""

Without a second thought, Doug leapt out of his chair

and said, **""Do you have a hat you could possibly spare?""**
","Yo, a neighbor was out there chillin' on his lawn",0
post,3jyjvk,2qh72,jokes,false,1441622769,https://old.reddit.com/r/Jokes/comments/3jyjvk/quick_oneliner_joke_why_are_pretty_women_like/,self.jokes,,"Because when they're not upright, they're grand! ",(Quick one-liner joke:) Why are pretty women like pianos?,3
post,3jyjfr,2qh72,jokes,false,1441622404,https://old.reddit.com/r/Jokes/comments/3jyjfr/how_can_you_tell_if_she_is_virgin_or_not/,self.jokes,,"Paddy was planning to get married and asked his doctor how he could tell if his bride is a virgin.

The doctor said, “Well, you need three things from a do it yourself shop. A can of red paint, a can of blue paint… and a shovel.”

Paddy asked, “And what do I do with these, doc?”

The doctor replied, “Before the wedding night, you paint one of your testicles red and the other one blue. If she says, ‘That’s the strangest pair of balls I ever saw.’, you hit her with the shovel.”
",How can you tell if she is virgin or not?,228
post,3jyj0q,2qh72,jokes,false,1441622059,https://old.reddit.com/r/Jokes/comments/3jyj0q/why_did_the_stop_sign_get_an_std/,self.jokes,,Because it had a 4-way.,Why did the stop sign get an STD?,0
post,3jyip5,2qh72,jokes,false,1441621812,https://old.reddit.com/r/Jokes/comments/3jyip5/guests/,self.jokes,,"There are two types of guests: the ones, who want to stay longer, and the ones, who want to go home asap. Strangely enough, these two types are normally found in married couples.

Read more at http://www.funny-jokes-quotes.com/daily-life-situations.html#UQbK0SvD6QcItByk.99",Guests,0
post,3jyid8,2qh72,jokes,false,1441621533,https://old.reddit.com/r/Jokes/comments/3jyid8/im_a_role_model/,self.jokes,,[deleted],I'm a role model!,1
post,3jyi34,2qh72,jokes,false,1441621298,https://old.reddit.com/r/Jokes/comments/3jyi34/a_computer_once_beat_me_at_chess/,self.jokes,,"It was no match for me at kick-boxing.







^shamelessly ^stolen ^from ^/u/enlighteningbug ^here: ^https://www.reddit.com/r/AskReddit/comments/3jul1x/what_critically_aclaimed_videogame_did_you_hate/cuslgfe",A computer once beat me at chess...,3
post,3jyhsg,2qh72,jokes,false,1441621041,https://old.reddit.com/r/Jokes/comments/3jyhsg/nsfwafter_a_round_of_golf/,self.jokes,,"a guy heads back to the club house. There, he sees a beautiful, blonde, big breasted woman, and naturally, he heads over to flirt with her. They hit it off, and decide to play a round together.

He is doing his best to impress, but she cleans his clock, winning by 9 strokes. Embarrassed, his manhood in question, she can tell he is hurt. But, she thinks he's sexy, so she suggests they go to the parking lot for a good ol' hummer in the backseat of his car. Needless to say, he enjoys himself and asks her to play golf tomorrow! 

She accepts, and every day that week, they play, she wins by a large amount, and afterwords he gets a BJ in his car. Though quite happy with the way things are going, he decides that he wants to seal the deal, and he invites her to his place for a romantic Saturday night dinner.

She shows up dressed to the 9s, the candles are lit, the steak is ready. They sit down to eat and a moment before his first bite she abruptly drops her silverware and exclaims, ""I can't do this anymore! I have to tell you something!""

Trying to comfort her, he says ""Of course, you can tell me anything! I'm sure it will be ok!"" To which she replies, ""I'm actually a MAN!""

His anger burns hotter than the sun, and he screams back, ""God damn you! You've been hitting off the women's tee all week!""

",[NSFW]After a round of golf...,892
post,3jyhgo,2qh72,jokes,false,1441620781,https://old.reddit.com/r/Jokes/comments/3jyhgo/why_are_asians_better_at_math_than_others/,self.jokes,,[deleted],Why are Asians better at math than others?,0
post,3jygis,2qh72,jokes,false,1441620039,https://old.reddit.com/r/Jokes/comments/3jygis/a_joke_for_blondes/,self.jokes,,"English is not my language but I hope I'll get it right.
So, it's the 1st intelligence championship for blondes. The stadium is packed with enthusiastic blondes and the runner up who has eliminated all other blonde contestants is ready for the question that will win her the title. The question is: what is the sum of 5 + 8. The countdown starts and we can see she is really struggling and at the end answers 12. The host goes all ""Oh, no, that was so close"" but the whole stadium starts chanting ""give her one more chance"". So they do give her one more chance. The question is: what is the sum of 5 + 7. Again, she struggles and at the end answers 13. The host goes all ""oh, no, that was so close"" but the whole stadium again starts chanting ""give her one more chance"". So they do. The question this time is: what is the sum of 5 + 5. She is really struggling and finally answers 10. The host goes ""yes, you did it"" and the whole stadium chants ""give her one more chance"".",A joke for blondes,2
post,3jyggb,2qh72,jokes,false,1441619993,https://old.reddit.com/r/Jokes/comments/3jyggb/the_trains_are_always_late/,self.jokes,,"A man was complaining to a railroad engineer. 
What's the use of having a train schedule if the trains are always late. 
The railroad engineer replied. 
How would we know they were late, if we didn't have a schedule? ",The Trains Are Always Late,3
post,3jyg8f,2qh72,jokes,false,1441619819,https://old.reddit.com/r/Jokes/comments/3jyg8f/my_mom_made_some_french_fries_for_you_guys/,self.jokes,,but you were dicks about it because they were potato quality.,My mom made some french fries for you guys...,3
post,3jyfda,2qh72,jokes,false,1441619112,https://old.reddit.com/r/Jokes/comments/3jyfda/sailors_and_lighters/,self.jokes,,"I was underway in the Pacific once when I witnessed one of my shipmates, up late, frantically attempting to smoke a cigarette. A burly Chief walks on-deck, roving as part of his duties - he didn't smoke himself.

One of the sailors asked the Chief if he had a Cigarette Lighter.

""Sure,"" the Chief said, ""Can I get a cigarette?""

Surprised, one of the junior sailors offered one to him. The Chief snatched it from his hand, and tossed it to the breeze - the stogie trailing with the wind into the ocean below.

""What was that all about, Chief?"" the younger sailor replied.

""I made the whole ship a cigarette lighter,"" he said, turning around and leaving.",Sailors and Lighters,1
post,3jyet8,2qh72,jokes,false,1441618659,https://old.reddit.com/r/Jokes/comments/3jyet8/first_experience_after_marriage/,self.jokes,,"A Delhi mother was lucky enough to see her 3 daughters get married the same year, so she called them after the wedding and told them

“Dont forget to text me your first night experience and text it in code”

So……. after a week, the 1st daughter texted

“NESCAFE”

and the next week the 2nd daughter text

“WILLS”

the mother being an intelligent woman went to get a Nescafe tin and read the label

“fantastic till the last drop”

went to her husband’s pack of WILLS cigarette and read
“Extra long, king size”

she smiled and said “not bad for their ages”.

After the next week, the 3rd daughter texted

“Indigo Delhi Hyderabad”,

the mother then called Indigo airways helpdesk to enquire about their Delhi Hyderabad flight and they replied

“it’s 5times daily, 7days a week, both ways and the flight duration is 75mins”.

Mother fainted",First Experience after marriage,1258
post,3jyeqc,2qh72,jokes,false,1441618593,https://old.reddit.com/r/Jokes/comments/3jyeqc/whats_the_difference_between_peanut_butter_and_jam/,self.jokes,,You can't peanut butter your dick into someone's ass.,What's the difference between peanut butter and jam.,0
post,3jydz3,2qh72,jokes,false,1441618004,https://old.reddit.com/r/Jokes/comments/3jydz3/parrot_with_no_legs/,self.jokes,,"A man suspected that his wife was cheating on him, but he could not find time to prove it since they worked opposite shifts. He soon came up with the idea to get a talking Parrot and hide it in the closet of the bedroom while he was gone.

He went to the local pet store and the clerk said ""we only have one Parrot that can talk real good, but he is sort of handicapped."" The husband asked, ""what's wrong with him?"" The clerk then told the man that the bird was born with no legs, so he holds himself up on the Perch by wrapping his long dick around it. The man agreed to buy the Parrot anyway.

Once the man arrived home, he put the Parrot in the bedroom closet and instructed the Parrot on what to do. Leaving the closet door partially open for the Parrot to see the bedroom, the man then left for work.

Arriving home the next morning the man noticed his wife had already left for work. He quickely went inside and began asking the Parrot, ""what have you seen?"" The Parrot replied ""You are right, your wife is cheating on you!"" ""Go on"", said the man. ""About a half an hour after you left, your wife came into the bedroom with another man! "" said the Parrot. ""Go on"", said the man. ""Then they took off all of their clothes and got onto the bed!"" ""Go on,""said the man. ""Then that guy started kissing your wife and sucking on her tits!"" said the Parrot. ""Then what happend?"", asked the man. ""Then that guy put his head between her legs and started licking her puss!"", said the Parrot. ""Then what?"" ,asked the man. ""I dont know"", said the Parrot, ""my dick got hard and I fell off the Perch!""




Couldn't find this anywhere after a brief scan - apologies if it's been posted before. Heard this as a young'un and it always tickled me",Parrot with no legs,59
post,3jycqc,2qh72,jokes,false,1441617003,https://old.reddit.com/r/Jokes/comments/3jycqc/heard_the_name_of_the_crappy_dollar_store_knock/,self.jokes,,[deleted],Heard the name of the crappy dollar store knock off of spitz sun flower seeds?,0
post,3jyb8m,2qh72,jokes,false,1441615818,https://old.reddit.com/r/Jokes/comments/3jyb8m/germany_are_welcoming_refugees_like_war_heroes/,self.jokes,,I'm mean.,Germany are welcoming refugees like war heroes because they had never had the chance to welcome the real thing.,0
post,3jyavg,2qh72,jokes,false,1441615521,https://old.reddit.com/r/Jokes/comments/3jyavg/2_elderly_couples_meet_up_one_afternoon/,self.jokes,,"The 2 husbands are chatting about what they've been up to recently. 
""We went to the most fantastic restaurant the other night"" says the first. 
""Which place was that?"" asks his friend. 
The first guy is really struggling to remember the name, and says ""Man, it's on the tip of my tongue, but I just can't remember.. What's the name of that flower, the one with sharp thorns on it, which is sometimes red or white, and has a nice smell?""

""Rose?"" Suggests the second. 

""Thats the one!!"" shouts the first, and then turns to his wife. 

""Rose!, what was the name of that restaurant we ate at the other night?"" 
",2 elderly couples meet up one afternoon,8
post,3jyap3,2qh72,jokes,false,1441615381,https://old.reddit.com/r/Jokes/comments/3jyap3/what_did_the_canadian_reddit_user_say/,self.jokes,,Ehhhhh lmao,What did the Canadian Reddit user say?,1
post,3jyacz,2qh72,jokes,false,1441615082,https://old.reddit.com/r/Jokes/comments/3jyacz/students_of_pathology_nsfw/,self.jokes,,"A professor in pathology is teaching his students what's important to become a good pathologist. In front of the group is a table with on it a dead body.  
""First of all,"" the professor says, ""It's important that you do not find anything disgusting.""  

To illustrate his point, the professors inserts his finger into the dead person's anus and subsequently puts his finger into his mouth. He then tells his students to do the same. Naturally there is some protest, but after a while all the students follow their teacher's example.  

When all the students have done this, the professor continues his lesson: ""Good. You have all proven that you do not find anything disgusting. Now for the second very important trait for a pathologist: eye to detail.   

Did anyone of you notice for example that I put my index finger into the dead person's anus, while it was my ring finger that I licked?""",Students of Pathology NSFW,171
post,3jy9l3,2qh72,jokes,false,1441614447,https://old.reddit.com/r/Jokes/comments/3jy9l3/what_did_the_alzheimers_patient_say_to_the_nurse/,self.jokes,,[deleted],What did the Alzheimer's patient say to the nurse?,0
post,3jy95b,2qh72,jokes,false,1441614092,https://old.reddit.com/r/Jokes/comments/3jy95b/are_my_testicles_black/,self.jokes,,"A man is in an accident and is placed on an oxygen mask to assist his breathing. 

His nurse checks on him and asks if there is anything he needs?

He say yes, could you check if my testicles are black?

She thinks, that is an odd request but decides to check for him as he looks very nervous.   

She looks at his testicles, flips them left and right and even rolls them in her hand to get a good look.  

After a few seconds she puts the sheet back down and notices the man smiling.  She says to him,""no sir your testicles are fine. Why are you smiling?""

He simply points at the mask, which she removes and he replies,""i just wanted to thank you for that experience, it was wonderful.   But, are my test results back?""",Are my testicles black?,310
post,3jy8tg,2qh72,jokes,false,1441613835,https://old.reddit.com/r/Jokes/comments/3jy8tg/there_was_a_guy_who_can_piss_real_limonade/,self.jokes,,"When it started to happen all his kids came up to him with cups, so he cam fill them with his lemonade, one of the kids had two cups,

""who's that for?"" The father asked

""It's for mommy, dad"" the kid replied.

""well, dont you worry about mommy, son, she will be drinking straight from the bottle"" - father",There was a guy who can piss real limonade,0
post,3jy8su,2qh72,jokes,false,1441613824,https://old.reddit.com/r/Jokes/comments/3jy8su/a_frenchman_an_englishman_and_a_russian_are/,self.jokes,,"The Frenchman says, “They must be French, they’re naked and they’re eating fruit.”

The Englishman replies with, “Clearly they’re English. Observe how politely the man is offering the woman the fruit.”

The Russian then notes, “They are Russian of course. They have nothing to wear, nothing to eat, and they think they are in paradise.”","A Frenchman, an Englishman and a Russian are admiring a painting of Adam and Eve in the garden of Eden...",72
post,3jy7ua,2qh72,jokes,false,1441613057,https://old.reddit.com/r/Jokes/comments/3jy7ua/eggs_and_toast_walk_into_a_bar/,self.jokes,,"And the bartender says, ""We don't serve breakfast here.""

",Eggs and Toast walk into a bar,1
post,3jy5ag,2qh72,jokes,false,1441611076,https://old.reddit.com/r/Jokes/comments/3jy5ag/how_did_the_farmer_find_the_sheep_in_the_tall/,self.jokes,,Satisfying.,How did the farmer find the sheep in the tall grass?,16
post,3jy4fz,2qh72,jokes,false,1441610425,https://old.reddit.com/r/Jokes/comments/3jy4fz/2_nuns_were_returning_to_the_monastery_after_a/,self.jokes,,"While they were crawling under the fence one nun turned to the other and said, ""I feel like a Marine!"" The other nun replied, ""Yeah, I do too. But where are we going to find one at this time of night?""",2 nuns were returning to the monastery after a night of drinking and partying in the town.,12
post,3jy3e3,2qh72,jokes,false,1441609654,https://old.reddit.com/r/Jokes/comments/3jy3e3/how_many_black_people_does_it_take_to_start_a_riot/,self.jokes,,-1,How many black people does it take to start a riot?,21
post,3jy39r,2qh72,jokes,false,1441609568,https://old.reddit.com/r/Jokes/comments/3jy39r/50_shades_of_hay/,self.jokes,,[50 shades of hay](http://imgur.com/YRGs7P0),50 shades of hay,0
post,3jy1vr,2qh72,jokes,false,1441608559,https://old.reddit.com/r/Jokes/comments/3jy1vr/an_irishman_walks_out_of_a_pub/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jy1vr/an_irishman_walks_out_of_a_pub/,,An Irishman walks out of a pub...,0
post,3jy16z,2qh72,jokes,false,1441608083,https://old.reddit.com/r/Jokes/comments/3jy16z/at_what_age_did_hitlers_uncle_try_to_molest_him_at/,self.jokes,,When he was nein.,At what age did Hitler's uncle try to molest him at?,0
post,3jy0xg,2qh72,jokes,false,1441607892,https://old.reddit.com/r/Jokes/comments/3jy0xg/why_does_crack_disproportionately_affect/,self.jokes,,[deleted],Why does crack disproportionately affect minorities?,0
post,3jxz7l,2qh72,jokes,false,1441606821,https://old.reddit.com/r/Jokes/comments/3jxz7l/i_was_in_a_restaurant_the_other_day/,self.jokes,,"I was in a restaurant the other day when suddenly I realized I desperately needed to pass gas. The music was really loud so i timed my gas with the beat of the music. After a couple of songs i started to feel better. I finished my coffee and noticed everyone was staring at me....
Then suddenly I remembered that I was listening to my ipod.",I was in a restaurant the other day...,3
post,3jxyet,2qh72,jokes,false,1441606239,https://old.reddit.com/r/Jokes/comments/3jxyet/whats_the_difference_between_a_chickpea_and_a/,self.jokes,,I've never paid to have a garbanzo bean on my chest ,Whats the difference between a chickpea and a garbanzo bean?,33
post,3jxydf,2qh72,jokes,false,1441606212,https://old.reddit.com/r/Jokes/comments/3jxydf/i_encountered_a_courteous_safe_driver_in_a/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jxydf/i_encountered_a_courteous_safe_driver_in_a/,,"I encountered a courteous, safe driver in a practical vehicle that had a marine corps decal on the rear windshield.",8
post,3jxyd4,2qh72,jokes,false,1441606204,https://old.reddit.com/r/Jokes/comments/3jxyd4/what_3_candies_do_you_find_in_school/,self.jokes,,"Redhots, DumDums, and smarties.",What 3 candies do you find in school?,1
post,3jxy2r,2qh72,jokes,false,1441605980,https://old.reddit.com/r/Jokes/comments/3jxy2r/if_you_guys_wanna_download_videos_of_your/,self.jokes,,[removed],If you guys wanna download videos of your favorite jokes on youtube then learn how to with this video.,1
post,3jxxz5,2qh72,jokes,false,1441605906,https://old.reddit.com/r/Jokes/comments/3jxxz5/girls_are_like_blackjack/,self.jokes,,I’m trying to go for 21 but I always hit on 14.,Girls are like blackjack.,115
post,3jxxbu,2qh72,jokes,false,1441605434,https://old.reddit.com/r/Jokes/comments/3jxxbu/today_is_labor_day/,self.jokes,,[deleted],Today is labor day!,0
post,3jxx9x,2qh72,jokes,false,1441605389,https://old.reddit.com/r/Jokes/comments/3jxx9x/do_you_know_what_i_am_looking_forward_to/,self.jokes,,[deleted],Do you know what I am looking forward to?,2
post,3jxw3m,2qh72,jokes,false,1441604628,https://old.reddit.com/r/Jokes/comments/3jxw3m/a_scotsman_stumbles_out_of_a_bar/,self.jokes,,"...completely wasted.  He was having trouble keeping his balance and knew he wouldn't make it walking home, so he found a nearby tree and propped himself up against it and proceeded to sleep it off.  A few minutes later, a couple of young lasses happen by.  They stop, and one looks at the other and says, ""Oh now, Mary, would you look at that?""

""What is it, June?""

""I've always wondered what was underneath a Scotsman's kilt!""

""Well have a look!""

So June bends over, lifts up the Scotsman's kilt and sees his penis there all in it's naked glory, and is pleasantly surprised.  ""Oh my, Mary,"" she exclaims.  ""Would you look at that!  It's beautiful!""

""Aye,"" says Mary.  ""You should leave him a present!""

So June thinks for a moment and gets an idea.  She takes the blue ribbon from her hair, ties it into a little bow around the Scotsman's penis, pulls the kilt down, and then she and Mary leave.

A few hours later, the Scotsman wakes up from his drunken slumber and has to take a piss.  So he goes around behind the tree, lifts up his kilt, and then he sees the blue ribbon.  Completely confused, he scratches his head for a moment and then exclaims, ""WELL, LADDEH!!  I DON' KNOW WHAR YA BE'N, BUT I'M GLAHD YA TOOK FARST PLACE!""",A Scotsman stumbles out of a bar...,9
post,3jxvn8,2qh72,jokes,false,1441604300,https://old.reddit.com/r/Jokes/comments/3jxvn8/9_out_of_10_people_enjoy_gang_rape/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jxvn8/9_out_of_10_people_enjoy_gang_rape/,,9 out of 10 people enjoy gang rape,6
post,3jxva0,2qh72,jokes,false,1441604066,https://old.reddit.com/r/Jokes/comments/3jxva0/you_know_why_i_wrap_duct_tape_around_my_hamsters/,self.jokes,,[deleted],You know why I wrap duct tape around my hamster's belly?,0
post,3jxv65,2qh72,jokes,false,1441603995,https://old.reddit.com/r/Jokes/comments/3jxv65/how_often_did_princess_sluttyness_get_laid/,self.jokes,,[deleted],How often did Princess Sluttyness get laid?,0
post,3jxv64,2qh72,jokes,false,1441603993,https://old.reddit.com/r/Jokes/comments/3jxv64/what_do_you_call_an_all_guy_christian_party/,self.jokes,,A suseJ fest,What do you call an all guy Christian party?,0
post,3jxuzi,2qh72,jokes,false,1441603868,https://old.reddit.com/r/Jokes/comments/3jxuzi/what_did_mick_jagger_say_when_he_walked_in_on/,self.jokes,,[removed],What did Mick Jagger say when he walked in on Hugh Hefner in bed with Dennis Weaver?,1
post,3jxuuo,2qh72,jokes,false,1441603790,https://old.reddit.com/r/Jokes/comments/3jxuuo/a_man_walks_into_a_bar/,self.jokes,,"he got a beer, waited the responsible 1 hour, and drove home.",A man walks into a bar..,0
post,3jxuhd,2qh72,jokes,false,1441603564,https://old.reddit.com/r/Jokes/comments/3jxuhd/a_wife_tells_her_husband_that_she_can_make_him/,self.jokes,,"The husband is baffled, ""Wha what? how is that even possible?""

The wife replies ""Well. you have the biggest dick of all your friends.""","A wife tells her husband that she can make him ""happy and sad"" at the same time.",89
post,3jxugb,2qh72,jokes,false,1441603551,https://old.reddit.com/r/Jokes/comments/3jxugb/early_christians_supported_marijuana_usage/,self.jokes,,Just think about how many get stoned.,Early christians supported marijuana usage.,3
post,3jxu9g,2qh72,jokes,false,1441603426,https://old.reddit.com/r/Jokes/comments/3jxu9g/an_irish_man_walks_out_of_a_bar/,self.jokes,,hahaha,An Irish man walks out of a bar,8
post,3jxu6x,2qh72,jokes,false,1441603381,https://old.reddit.com/r/Jokes/comments/3jxu6x/what_is_the_hardest_part_of_eating_a_vegetable/,self.jokes,,The wheelchair.,What is the hardest part of eating a vegetable?,3
post,3jxu62,2qh72,jokes,false,1441603368,https://old.reddit.com/r/Jokes/comments/3jxu62/how_do_you_make_a_giraffe_go_to_war/,self.jokes,,You Giraffed it,How do you make a Giraffe go to war?,2
post,3jxtre,2qh72,jokes,false,1441603132,https://old.reddit.com/r/Jokes/comments/3jxtre/what_do_you_call_a_half_elephant_half_rhinoceros/,self.jokes,,"An abomination.

","What do you call a half elephant, half rhinoceros?",0
post,3jxt8i,2qh72,jokes,false,1441602789,https://old.reddit.com/r/Jokes/comments/3jxt8i/my_cute_kitten/,self.jokes,,"Aww, wrong sub.",My cute kitten,1
post,3jxt12,2qh72,jokes,false,1441602658,https://old.reddit.com/r/Jokes/comments/3jxt12/what_does_a_baby_in_a_blender_sound_like/,self.jokes,,"I don't know, I couldn't hear it over the sound of my masturbating.",What does a baby in a blender sound like?,0
post,3jxt0u,2qh72,jokes,false,1441602650,https://old.reddit.com/r/Jokes/comments/3jxt0u/what_did_mick_jagger_say_when_he_walked_in_on/,self.jokes,,[removed],What did Mick Jagger say when he walked in on Hugh Hefner having sex with Dennis Weaver?,1
post,3jxslq,2qh72,jokes,false,1441602383,https://old.reddit.com/r/Jokes/comments/3jxslq/a_man_walks_into_a_brothel/,self.jokes,,"He approaches the lady at the front desk and says, ""Hi, I would like to purchase some sex please."" 
The lady just smiled and replied, ""Ok, here is the board with the different priced women. All are currently available right now so choose whoever you'd like.""
The man looking a bit concerned said, ""Well you see, I only have $20. What will that do for me?""
""Oh...wellll I will just have to give you the cheapest lady then. But don't worry, you're not the first! Here is your room key and she'll be waiting for you in room D."" The lady replied. 
Excited and nervous the man ran to his room. After about 10 minutes he came out sprinting back to the front desk and frantically rang the bell repeatedly. The lady came out curious what he was so frantic about.
""Yes? What can I help you with?"" She asked.
The man exclaimed, ""I went in the room and noticed my girl was acting strange and not very responsive, but I disregarded it and started getting my thang on. Then all of a sudden puss started pouring out of her nose and mouth! We need to call an ambulance or something!""
The lady at the front desk just replies, ""Ohhh, don't worry about that. Hey Doug! The dead chick in room D is full again!"" ",A man walks into a brothel...,1
post,3jxsi7,2qh72,jokes,false,1441602315,https://old.reddit.com/r/Jokes/comments/3jxsi7/a_guy_walks_into_a_pub/,self.jokes,,he was hiding from the police after they shot his family for j walking,A guy walks into a pub,0
post,3jxqvl,2qh72,jokes,false,1441601297,https://old.reddit.com/r/Jokes/comments/3jxqvl/whats_worse_than_lobsters_on_your_piano/,self.jokes,,Syphilis,What's worse than lobsters on your piano?,3
post,3jxqcy,2qh72,jokes,false,1441601002,https://old.reddit.com/r/Jokes/comments/3jxqcy/a_guy_walks_into_a_pub/,self.jokes,,[deleted],A guy walks into a pub...,0
post,3jxq4h,2qh72,jokes,false,1441600860,https://old.reddit.com/r/Jokes/comments/3jxq4h/why_do_the_dutch_value_geometry_so_much/,self.jokes,,[deleted],Why do the Dutch value geometry so much?,4
post,3jxplf,2qh72,jokes,false,1441600536,https://old.reddit.com/r/Jokes/comments/3jxplf/my_girlfriend_keeps_thinking_iam_leaving_her/,self.jokes,,"She fell on the floor one day and took a hit, now whenever i bump the lid she's always saying goodbye. i think i need to get my laptop fixed.",My girlfriend keeps thinking iam leaving her...,0
post,3jxovn,2qh72,jokes,false,1441600127,https://old.reddit.com/r/Jokes/comments/3jxovn/two_men_are_at_dinner/,self.jokes,,"Two men are sitting at dinner one night, when one looks out the window and asks the other,""Which do you think is closer: the moon or Miami?""

The other man replies, ""Well... you can't SEE Miami.""",Two men are at dinner,0
post,3jxojb,2qh72,jokes,false,1441599898,https://old.reddit.com/r/Jokes/comments/3jxojb/what_are_the_consequences_of_smoking_weed/,self.jokes,,The reefercussions,What are the consequences of smoking weed?,2
post,3jxnf9,2qh72,jokes,false,1441599204,https://old.reddit.com/r/Jokes/comments/3jxnf9/three_men_have_to_share_a_bed/,self.jokes,,"They're on a ski trip together, and due to a clerical error there is only one room left in the lodge. There is only one large bed, and there are no cots.

So the three pile in and try to keep their distance.

The next morning they wake up, and the man sleeping on the left edge of the bed says:

""I had the best sleep! I dreamed that a beautiful Scandinavian goddess was making love to me, her lips were like pillows!""

The man sleeping at the right edge of the bed says ""So did I! I dreamed I was fucking a blonde bombshell!""
 He turns to the man in the middle and asks ""What did you dream about?"" 

He replies:

""Skiing.""",Three men have to share a bed,11
post,3jxmtg,2qh72,jokes,false,1441598848,https://old.reddit.com/r/Jokes/comments/3jxmtg/i_asked_my_heart/,self.jokes,,[deleted],I asked my Heart...,0
post,3jxmsg,2qh72,jokes,false,1441598829,https://old.reddit.com/r/Jokes/comments/3jxmsg/i_think_my_neighbor_is_stalking_me/,self.jokes,,as I saw her googling my name on her computer last night.I saw it through my telescope.,I think my neighbor is stalking me...,3
post,3jxmqj,2qh72,jokes,false,1441598802,https://old.reddit.com/r/Jokes/comments/3jxmqj/a_young_mans_grandfather_dies/,self.jokes,,"He asks his Grandmother how he died.

She said "" Well every Sunday We would make love to the sound of the church bells, they were slow enough for us.""

The young man asked ""But how did he die then?""

She replied "" He would still be alive if it wasn't for that damn Ice Cream truck.""",A young man's Grandfather dies.,7
post,3jxmqf,2qh72,jokes,false,1441598801,https://old.reddit.com/r/Jokes/comments/3jxmqf/two_guys_walk_into_a_dinner/,self.jokes,,"They sit down and the waitress takes their order.
   ""Two cheese burgers and fries.""
They watch as she walks to the kitchen window and gives the cook the order slip. The cook reads it and turns to the cooler and grabs a hand full of ground beef. He sticks it in his arm pit and brings his arm down smashing it flat, then tosses it on the grill. They watch again in disbelief as he grabs another hand full of ground beef and again sticks it in his arm pit and smashes it flat with his big sweaty arm, then drops in down beside the other one.
    They call the waitress over and ask her what the hell is he doing preparing food like that and she replies, ""Oh that's nothing you should be here when he pokes the poles in the doughnuts.""",Two guys walk into a dinner,9
post,3jxmju,2qh72,jokes,false,1441598706,https://old.reddit.com/r/Jokes/comments/3jxmju/an_irish_man_walks_into_a_bar/,self.jokes,,.,An Irish man walks into a bar.,0
post,3jxklb,2qh72,jokes,false,1441597576,https://old.reddit.com/r/Jokes/comments/3jxklb/how_do_you_get_a_jewish_girls_number/,self.jokes,,you ask her to roll her sleeves up.,How do you get a Jewish girls number?,1
post,3jxkjn,2qh72,jokes,false,1441597550,https://old.reddit.com/r/Jokes/comments/3jxkjn/why_should_you_never_take_a_pig_out_on_a_date/,self.jokes,,She might squeal on you.,Why should you never take a pig out on a date?,7
post,3jxka4,2qh72,jokes,false,1441597390,https://old.reddit.com/r/Jokes/comments/3jxka4/two_jews_walk_by_a_christian_church/,self.jokes,,"There is a sign on the door that says, ""convert to Christianity and receive $100"". One of them speaks up and says, ""I'm going in."" His friend says ""you're really going to change religions for $100?"" 
""A $100 is a $100, I'm doing it!"" And he walks inside. 
A few minutes later he walks back out and his friend says, ""Well? Did you get the money?""
He replies, ""Oh, that's all you people think about isn't it?""
",Two Jews walk by a Christian church. . .,31
post,3jxjj2,2qh72,jokes,false,1441596948,https://old.reddit.com/r/Jokes/comments/3jxjj2/what_did_the_forward_rooster_say/,self.jokes,,Cock a doodle do. What did the backward rooster say? Doodle doodle cock. WHAT did the gay rooster say? Any cock will do.,What did the forward rooster say?,2
post,3jxj43,2qh72,jokes,false,1441596716,https://old.reddit.com/r/Jokes/comments/3jxj43/on_his_20th_wedding_anniversary_a_man_proposes_a/,self.jokes,,"He's surprised when she slaps him across the face. ""What was that for?"" he asks. 

""For 20 years of bad sex.""

The man then slaps his wife across the face. ""What was that for?"" she demands.

""For knowing the difference.""
","On his 20th wedding anniversary, a man proposes a toast to his wife.",3
post,3jxipj,2qh72,jokes,false,1441596521,https://old.reddit.com/r/Jokes/comments/3jxipj/whats_the_difference_between_a_porsche_and_a_pile/,self.jokes,,"When I see a porsche on the street I think ""hey, thats a nice car,"" but when I see a pile of dead babies, I scream, ""OH DEAR GOD WHY? WHY GOD WHY? WHERE IS THE MONSTER WHO DID THIS? NO GOD NOOO!",What's the difference between a porsche and a pile of dead babies?,0
post,3jxif8,2qh72,jokes,false,1441596359,https://old.reddit.com/r/Jokes/comments/3jxif8/the_lone_ranger/,self.jokes,,[deleted],The Lone Ranger...,1
post,3jxibi,2qh72,jokes,false,1441596305,https://old.reddit.com/r/Jokes/comments/3jxibi/whats_brown_and_sticky/,self.jokes,,A stick.,What's brown and sticky?,11
post,3jxhy3,2qh72,jokes,false,1441596091,https://old.reddit.com/r/Jokes/comments/3jxhy3/heaven/,self.jokes,,[deleted],Heaven,21
post,3jxhbr,2qh72,jokes,false,1441595751,https://old.reddit.com/r/Jokes/comments/3jxhbr/fuck_you/,self.jokes,,[removed],FUCK YOU,0
post,3jxgjc,2qh72,jokes,false,1441595285,https://old.reddit.com/r/Jokes/comments/3jxgjc/a_jew_a_catholic_and_a_colored_boy_go_to_heaven/,self.jokes,,"They get to the pearly gates and are surrounded by clocks.  So the Jew asks St. Peter "" Yo Pete what's up with all these clocks?""  St. Peter looks over his tri focal glasses and says"" Every time you masturbate the clock goes around once, yours is right over there.  It goes around about once a week.""  The catholic giggles a little and the Jew asks "" where is his?"" pointing to the catholic.  "" His is right over there, goes around once a day and twice on Sunday."" St Peter says with a smirk.  The Jew and the catholic look at the colored boy whose eyes are as big as saucers with a horrified look on his face.  "" What about him?""  ""Oh his in Jesus's  room, he uses it for a fan.  ","A Jew, a Catholic and a Colored boy go to heaven.",4
post,3jxg1z,2qh72,jokes,false,1441595009,https://old.reddit.com/r/Jokes/comments/3jxg1z/some_pages_troll_us_by_making_a_pixel_or_two_on/,self.jokes,,I just can't put my finger on it.,Some pages troll us by making a pixel or two on the page black so that we think it's a smudge... why would anyone do that?,2
post,3jxfn7,2qh72,jokes,false,1441594780,https://old.reddit.com/r/Jokes/comments/3jxfn7/poor_jimmy_was_being_teased_by_two_of_his_friends/,self.jokes,,[deleted],Poor Jimmy was being teased by two of his friends...,0
post,3jxeyx,2qh72,jokes,false,1441594376,https://old.reddit.com/r/Jokes/comments/3jxeyx/im_going_to_the_bathroom_to_take_a_dump/,self.jokes,,Can I get you anything?,I'm going to the bathroom to take a dump,0
post,3jxece,2qh72,jokes,false,1441594044,https://old.reddit.com/r/Jokes/comments/3jxece/whats_the_difference_between_an_oyster_fisherman/,self.jokes,,The oyster fisherman shucks between fits.,What's the difference between an oyster fisherman with epilepsy and a prostitute with diarrhea?,94
post,3jxdv8,2qh72,jokes,false,1441593751,https://old.reddit.com/r/Jokes/comments/3jxdv8/jazz_clubs/,self.jokes,,"My friend was telling me about how much he loves jazz music, and he was telling me about a jazz club he goes to.

I also go to a jazz club, called ""Hot Jazz in Your Face"", and I made my friend aware of this.

He asked, ""Where can I find it?""

I replied, ""Oh, they closed it down...""

""Why did they close it?""

""People just stopped... coming...""",Jazz Clubs,0
post,3jxdh8,2qh72,jokes,false,1441593524,https://old.reddit.com/r/Jokes/comments/3jxdh8/i_went_to_the_pub_the_other_night/,self.jokes,,"I went to the pub the other night.  There were three rather hefty ladies having a rowdy good time.  Their accent appeared to be Scottish so I approached and asked, ""Hello ladies, are you three lassies from Scotland?""  One of them angrily screeched, ""It's Wales you bloody idiot, Wales!""  So I apologized and replied, ""I'm terribly sorry.  Are you three whales from Scotland?""

PS: Probably an oldie but I just heard it recently.",I went to the pub the other night,16
post,3jxda2,2qh72,jokes,false,1441593417,https://old.reddit.com/r/Jokes/comments/3jxda2/a_guy_in_a_jeep_stops_to_put_air_in_his_tire_at_a/,self.jokes,,The air costs 25 cents.  He walks into the gas station and hands the attendant 25 cents.  The attendant looks at his jeep with a New England Patriots cover on the spare tire and says here you can have your quarterback.,A guy in a jeep stops to put air in his tire at a gas station.,3
post,3jxcxb,2qh72,jokes,false,1441593229,https://old.reddit.com/r/Jokes/comments/3jxcxb/a_family_walks_into_a_hotel/,self.jokes,,[deleted],A family walks into a hotel...,1
post,3jxcht,2qh72,jokes,false,1441593022,https://old.reddit.com/r/Jokes/comments/3jxcht/how_do_you_bury_a_pothead/,self.jokes,,Coughin',How do you bury a pothead?,3
post,3jxcb7,2qh72,jokes,false,1441592920,https://old.reddit.com/r/Jokes/comments/3jxcb7/a_tactile_reply_in_tense_situations/,self.jokes,,"Once asked, ""What is a solid reply to a strong, hearty 'Fuck You'?"" the editor of Playboy blithely remarked, ""Fuck yourself. You'll get more pussy that way."" 

A non traditional joke. Stay out trouble this weekend!",A tactile reply in tense situations,3
post,3jxc9o,2qh72,jokes,false,1441592889,https://old.reddit.com/r/Jokes/comments/3jxc9o/what_do_you_do_when_your_dishwasher_stops_working/,self.jokes,,"Beat it until she starts again.
",What do you do when your dishwasher stops working?,0
post,3jxc02,2qh72,jokes,false,1441592728,https://old.reddit.com/r/Jokes/comments/3jxc02/apparently_trump_wants_to_outlaw_preshredded/,self.jokes,,...he keeps going on and on about how he wants to make America grate again...,Apparently Trump wants to outlaw pre-shredded cheese...,39
post,3jxasl,2qh72,jokes,false,1441592064,https://old.reddit.com/r/Jokes/comments/3jxasl/what_does_korean_food_taste_like/,self.jokes,,Chinese food.,What does Korean food taste like?,0
post,3jx9zf,2qh72,jokes,false,1441591616,https://old.reddit.com/r/Jokes/comments/3jx9zf/my_favorite_pokemon_is_electrode/,self.jokes,,[deleted],My favorite Pokemon is Electrode.,1
post,3jx8zw,2qh72,jokes,false,1441591106,https://old.reddit.com/r/Jokes/comments/3jx8zw/a_dog_is_walking_through_the_forest/,self.jokes,,"...and runs into his old friend , an owl. ""It's been a long time, how's it going?"" the dog inquires. ""Great, life's a hoot,"" replies the owl, ""how are you?""  ""For me, it's been ruff.""",A dog is walking through the forest...,0
post,3jx73q,2qh72,jokes,false,1441590098,https://old.reddit.com/r/Jokes/comments/3jx73q/i_ate_a_stary_poprock_that_stuck_to_my_palm/,self.jokes,,[deleted],I ate a stary poprock that stuck to my palm...,1
post,3jx6x3,2qh72,jokes,false,1441590001,https://old.reddit.com/r/Jokes/comments/3jx6x3/whats_the_difference_between_a_canoe_and_a_jewish/,self.jokes,,[deleted],What's the difference between a canoe and a Jewish person?,1
post,3jx6vl,2qh72,jokes,false,1441589978,https://old.reddit.com/r/Jokes/comments/3jx6vl/dont_take_life_too_seriously/,self.jokes,,[deleted],Don't take life too seriously,5
post,3jx6pk,2qh72,jokes,false,1441589899,https://old.reddit.com/r/Jokes/comments/3jx6pk/chris_hanson_dressing_up_as_arnold_schwarzenegger/,self.jokes,,[deleted],Chris Hanson dressing up as Arnold Schwarzenegger....,0
post,3jx6du,2qh72,jokes,false,1441589741,https://old.reddit.com/r/Jokes/comments/3jx6du/kaliningrad/,self.jokes,,[deleted],Kaliningrad,1
post,3jx6db,2qh72,jokes,false,1441589733,https://old.reddit.com/r/Jokes/comments/3jx6db/i_was_on_this_plane_once/,self.jokes,,"I was on this plane once. And I'm sittin' there and the captain comes on and he does his whole, ""We'll be cruising at 35,000 feet,"" then he puts the mike down but he forgets to turn it off. Then he turns to the copilot and goes, ""You know, all I could go for right now is a blow job and a cup of coffee."" So the stewardess goes bombin' up from the back of the plane to tell him the mic's still on, and this guy behind me goes, ""Hey hon, don't forget the coffee!""

From Good Will Hunting",I was on this plane once,4
post,3jx5um,2qh72,jokes,false,1441589460,https://old.reddit.com/r/Jokes/comments/3jx5um/three_oaps_are_sitting_in_a_retirement_home/,self.jokes,,[removed],Three OAP's are sitting in a retirement home discussing life,1
post,3jx5fj,2qh72,jokes,false,1441589245,https://old.reddit.com/r/Jokes/comments/3jx5fj/why_do_scotsmen_wear_kilts/,self.jokes,,[deleted],Why do Scotsmen wear kilts?,1
post,3jx5cl,2qh72,jokes,false,1441589197,https://old.reddit.com/r/Jokes/comments/3jx5cl/my_wife_wants_to_have_the_baby_listen_to/,self.jokes,,Would an ipod nano or shuffle be easier to get up there?,My wife wants to have the baby listen to classical music while in the womb.,21
post,3jx533,2qh72,jokes,false,1441589065,https://old.reddit.com/r/Jokes/comments/3jx533/what_do_you_call_a_multiple_choice_dad_joke/,self.jokes,,A pop quiz.,What do you call a multiple choice dad joke?,2
post,3jx47h,2qh72,jokes,false,1441588610,https://old.reddit.com/r/Jokes/comments/3jx47h/how_do_you_make_five_pounds_of_fat_look_good/,self.jokes,,[deleted],How do you make five pounds of fat look good?,3
post,3jx3vz,2qh72,jokes,false,1441588432,https://old.reddit.com/r/Jokes/comments/3jx3vz/salesman/,self.jokes,," A sales company has particular trouble selling bibles. One day, a man comes in with a job application and says, ""l-l-l-l'd l-l-l-l-l-like t-t-t-t-t-to b-b-b-b- b-be a b-b-b-bible salesman, s-s-s-sir."" lnititally, he doesn't want to give the job to this man, but decided to try him out.

After three weeks, the manager is looking at the charts and realizes that the newest guy is selling the most copies. Amazed, he calls him in to his office. ""You've only worked here for three weeks and you've already sold more copies than anyone else here! How do you do it?""

""W-w-w-w-w-well, l g-g-g-go up t-t-t-t-to th-the d-d-d-door and-d-d l-l--l s-s-s-say, w-w-w-w-would y-y-y-y-y-y-you l-l-l-l-l-like t-t-to b-b-b-b-buy a  b-b-b-bible, or w-w-w-would y-y-you l-l-l-like m-m-me t-t-t-to r-r-r-r-read it t-t-t-t-t-to y-y-y-you?"" ",Salesman,62
post,3jx352,2qh72,jokes,false,1441588008,https://old.reddit.com/r/Jokes/comments/3jx352/your_mother_has_the_prettiest_teeth_i_ever_came/,self.jokes,,Your mother has the prettiest teeth I ever came across.,Your mother has the prettiest teeth I ever came across.,17
post,3jx2dz,2qh72,jokes,false,1441587619,https://old.reddit.com/r/Jokes/comments/3jx2dz/what_did_the_buffalo_say_to_his_son_when_he_left/,self.jokes,,[deleted],What did the buffalo say to his son when he left for college?,50
post,3jx28u,2qh72,jokes,false,1441587549,https://old.reddit.com/r/Jokes/comments/3jx28u/whats_more_awkward_than_walking_in_on_your/,self.jokes,,[deleted],What's more awkward than walking in on your parents having sex?,0
post,3jx1y1,2qh72,jokes,false,1441587384,https://old.reddit.com/r/Jokes/comments/3jx1y1/whats_the_strongest_muscle_on_a_pig/,self.jokes,,The hamstring.,What's the strongest muscle on a pig?,4
post,3jx1lt,2qh72,jokes,false,1441587193,https://old.reddit.com/r/Jokes/comments/3jx1lt/brotherly_love/,self.jokes,,"A new Irish pub opens in downtown New York. On the first day, an Irishman walks in and orders three pints of Guinness.


He takes a sip from the first one, then a sip from the second and finally a sip from the third. He does this in turn until all pints are empty. This goes on every day for a few weeks, and since the barkeeper has never seen anything like this, he asks about this peculiar drinking habit one day:


“See”, the Irishman says, “I used to go for a pint together with my two brothers. But Paddy, my older brother, moved back home to Kerry and my younger brother, Sean, moved to Boston. So, now that it’s just me, I order a pint for each of them as well. We agreed as long we’re all still drawing breath, we’ll raise a glass together, just like we used to. Sláinte!”


Thinking this is a lovely tradition, the barman continues to serve his patron three pints and watches him drink them sip by sip every evening for the next few months. One day, however, the man comes in and orders *just two pints*. He takes turns drinking them as usual and goes home. This goes on for a few days, before the barkeeper works up the courage to talk to him:


“You told me about your tradition, that as long as the three of you were still alive, you’d continue drinking together. I am so sorry to hear about your brother passing. Drinks are on the house today.”


To which the Irishman responds.


“Cheers, but both my brothers are doing fine. It’s just my doctor has prescribed me a new type of medicine and told me that *I* need to stop drinking.”
",Brotherly Love,34
post,3jx0je,2qh72,jokes,false,1441586594,https://old.reddit.com/r/Jokes/comments/3jx0je/a_man_who_thinks_his_wife_might_be_cheating_on/,self.jokes,,"...The hit-man says it will cost $5000. The man says that's fine but he wants to watch. The hit-man agrees so they find a spot on a nearby roof and wait for the wife to get home. 

Eventually the wife comes home and she's with a guy.
The husband is furious but still not sure if she is cheating yet so they wait some more.

Eventually the hit-man pulls out his binoculars and after about 30 seconds he says ""oh ya she's cheating on you. What do you want me to do?"".

The irate husband says ""Put a bullet in her head and while you're at it put a bullet in the guys dick as well"".

The hitman replies ""Ok, but that's going to cost you another $5000. The good news is I'm only going to need one bullet."" ",A man who thinks his wife might be cheating on him hires a hit-man..,154
post,3jx029,2qh72,jokes,false,1441586358,https://old.reddit.com/r/Jokes/comments/3jx029/you_know_what_they_say_about_moldy_tents/,self.jokes,,That mold is intense. ,You know what they say about moldy tents....,4
post,3jwyjt,2qh72,jokes,false,1441585657,https://old.reddit.com/r/Jokes/comments/3jwyjt/knock_knock/,self.jokes,,"Who's there?

9/11.
9/11 who?
I though you'd never forget.",Knock Knock.,0
post,3jwxs8,2qh72,jokes,false,1441585246,https://old.reddit.com/r/Jokes/comments/3jwxs8/so_this_joke_is_only_half_finished/,self.jokes,,[deleted],So This Joke Is Only Half Finished...,0
post,3jwx1w,2qh72,jokes,false,1441584876,https://old.reddit.com/r/Jokes/comments/3jwx1w/hand_is_all_you_need/,self.jokes,,"Mark: I hope tonight will be a night to remember!

John: A hand is all you really need.

Mark: A hand is all I got.",Hand is all you need ...,0
post,3jwwx2,2qh72,jokes,false,1441584805,https://old.reddit.com/r/Jokes/comments/3jwwx2/whats_the_difference_between_a_duck_and_george/,self.jokes,,[deleted],What's the difference between a duck and George Washington?,0
post,3jwvmf,2qh72,jokes,false,1441584142,https://old.reddit.com/r/Jokes/comments/3jwvmf/hand_is_all_i_need/,self.jokes,,[deleted],Hand is all I need.,1
post,3jwvhj,2qh72,jokes,false,1441584074,https://old.reddit.com/r/Jokes/comments/3jwvhj/a_woman_is_late_to_a_fight_she_takes_a_seat_next/,self.jokes,,"""How many cocks have been beaten?"" she asks.

""None, until now,"" says a man with a smile.",A woman is late to a fight. She takes a seat next to several men.,0
post,3jwuul,2qh72,jokes,false,1441583754,https://old.reddit.com/r/Jokes/comments/3jwuul/a_man_goes_to_his_friend_for_advice_as_his_wife/,self.jokes,,"His friend tells him to go home looking angry, and take of his clothes and have a shower as that would help mask his breath and erase the smell.the man agrees and rides his bike home after having a few drinks, he goes home looking angry and takes off his clothes just when he's about to enter the bathroom, his wife asks him if he's drunk. He replies no, im just having a shower and the wife says why didn't you take off your helmet if you're having a shower. And the man dies...",A man goes to his friend for advice as his wife always finds out he's drunk when he comes home,0
post,3jwtzn,2qh72,jokes,false,1441583280,https://old.reddit.com/r/Jokes/comments/3jwtzn/what_is_the_blonde_doing_when_she_holds_her_hands/,self.jokes,,[deleted],What is the blonde doing when she holds her hands tightly over her ears?,2
post,3jwtso,2qh72,jokes,false,1441583195,https://old.reddit.com/r/Jokes/comments/3jwtso/so_jesus_walks_into_a_bar/,self.jokes,,[deleted],So Jesus walks into a bar...,0
post,3jwto7,2qh72,jokes,false,1441583132,https://old.reddit.com/r/Jokes/comments/3jwto7/a_line_from_my_grandfather/,self.jokes,,[deleted],A line from my grandfather,0
post,3jwsrq,2qh72,jokes,false,1441582618,https://old.reddit.com/r/Jokes/comments/3jwsrq/my_wife_asked_if_i_was_coming_to_our_daughters/,self.jokes,,"I was, but I paused the video, pulled up my pants, and denied it.",My wife asked if I was coming to our daughter's dance recital...,9
post,3jwskd,2qh72,jokes,false,1441582488,https://old.reddit.com/r/Jokes/comments/3jwskd/the_deli/,self.jokes,,"I was once arrested for scalping low numbers in the deli at the grocery. 


                      Note - There is a funny comedian, Steve Wright, he said this one on the tonight show back in the Carson days. He was funny as hell! ",The Deli,0
post,3jwsfv,2qh72,jokes,false,1441582420,https://old.reddit.com/r/Jokes/comments/3jwsfv/did_you_hear_about_the_blonde_actress_that/,self.jokes,,"Reese Witherspoon?

No with her fork!",Did you hear about the blonde actress that stabbed her husband with a fork? Reese something...,2
post,3jwrn9,2qh72,jokes,false,1441581992,https://old.reddit.com/r/Jokes/comments/3jwrn9/how_do_you_build_suspense/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jwrn9/how_do_you_build_suspense/,,How do you build suspense?,0
post,3jwrmh,2qh72,jokes,false,1441581981,https://old.reddit.com/r/Jokes/comments/3jwrmh/whats_a_convicted_criminal_who_plays_with_other/,self.jokes,,[deleted],What's a convicted criminal who plays with other people's emotions?,1
post,3jwrj3,2qh72,jokes,false,1441581928,https://old.reddit.com/r/Jokes/comments/3jwrj3/hey_girl_you_got_a_kind_face/,self.jokes,,[deleted],"Hey girl, you got a kind face....",0
post,3jwqs8,2qh72,jokes,false,1441581516,https://old.reddit.com/r/Jokes/comments/3jwqs8/where_on_earth_can_you_find_the_highest/,self.jokes,,In the atmosphere.,Where on Earth can you find the highest concentration of Jews?,1
post,3jwp7o,2qh72,jokes,false,1441580706,https://old.reddit.com/r/Jokes/comments/3jwp7o/an_elderly_woman_had_her_purse_stolen_by_a_man_in/,self.jokes,,"And as he wheeled away she yelled ""You can hide, but you can't run!""",An elderly woman had her purse stolen by a man in a wheelchair...,1
post,3jwp6a,2qh72,jokes,false,1441580680,https://old.reddit.com/r/Jokes/comments/3jwp6a/mr_president_another_two_brazilian_soldiers_were/,self.jokes,,[deleted],"""Mr. President, another two Brazilian soldiers were killed yesterday in Iraq.""",0
post,3jwor6,2qh72,jokes,false,1441580460,https://old.reddit.com/r/Jokes/comments/3jwor6/narcos_sushi_thought_for_the_day_how_have_i_never/,self.jokes,,That is all.  You may laugh now.,"Narcos + Sushi thought for the day: How have I never come across a roll called the ""Pablo Escolar""?",0
post,3jwo37,2qh72,jokes,false,1441580138,https://old.reddit.com/r/Jokes/comments/3jwo37/how_do_you_avoid_the_constant_apple_reboot_loop/,self.jokes,,Don’t make a third movie,How do you avoid the constant Apple reboot loop?,1
post,3jwo0g,2qh72,jokes,false,1441580095,https://old.reddit.com/r/Jokes/comments/3jwo0g/im_throwing_a_party_for_people_who_cant_ejaculate/,self.jokes,,Tell me if you can come.,I'm throwing a party for people who can't ejaculate...,0
post,3jwmn3,2qh72,jokes,false,1441579363,https://old.reddit.com/r/Jokes/comments/3jwmn3/how_many_psychiatrist_does_it_take_to_change_a/,self.jokes,,"Just one, but it takes a really long time, and the lightbulb has to want to change...",How many psychiatrist does it take to change a lightbulb?,5
post,3jwlxm,2qh72,jokes,false,1441579008,https://old.reddit.com/r/Jokes/comments/3jwlxm/a_guy_walks_into_a_pub/,self.jokes,,"...And sees a sign hanging over the bar that reads: CHEESEBURGER: $1.50 CHICKEN SANDWICH: $2.50 HAND JOB: $10.00 He walks up to the bar and beckons one of the three exceptionally attractive blondes serving drinks. ""Can I help you?"" she asks. ""I was wondering,"" whispers the man. ""Are you the one who gives the hand jobs?"" ""Yes,"" she purrs. ""I am."" The man replies, ""Well, wash your hands. I want a cheeseburger.""",A guy walks into a pub...,8814
post,3jwluq,2qh72,jokes,false,1441578962,https://old.reddit.com/r/Jokes/comments/3jwluq/lay_off/,self.jokes,,[deleted],Lay off!,1
post,3jwlsh,2qh72,jokes,false,1441578928,https://old.reddit.com/r/Jokes/comments/3jwlsh/your_mom_is_like_rambo/,self.jokes,,[deleted],Your mom is like rambo,0
post,3jwlhb,2qh72,jokes,false,1441578761,https://old.reddit.com/r/Jokes/comments/3jwlhb/what_is_another_name_for_a_goofy_stoner_grin/,self.jokes,,[deleted],What is another name for a goofy stoner grin?,0
post,3jwlf8,2qh72,jokes,false,1441578733,https://old.reddit.com/r/Jokes/comments/3jwlf8/happy_times_with_grandma/,self.jokes,,"One day I was eating my grandma out. 

Suddenly I tasted horse semen. 

""I thought"" Oh yeah, that's how she died. ",Happy times with grandma,0
post,3jwl9z,2qh72,jokes,false,1441578659,https://old.reddit.com/r/Jokes/comments/3jwl9z/what_do_you_get_when_you_sit_under_a_cow/,self.jokes,,A pat on the head. ,What do you get when you sit under a cow?,3
post,3jwl75,2qh72,jokes,false,1441578618,https://old.reddit.com/r/Jokes/comments/3jwl75/whats_worse_than_lobsters_on_your_piano/,self.jokes,,Crabs on your organ.  (still my favorite joke from grade school),What's worse than lobsters on your piano?,30
post,3jwl65,2qh72,jokes,false,1441578606,https://old.reddit.com/r/Jokes/comments/3jwl65/whats_the_difference_between_a_fish_and_a/,self.jokes,,Fish muck about in fountains…,What’s the difference between a fish and a mountain goat?,10
post,3jwjrl,2qh72,jokes,false,1441577881,https://old.reddit.com/r/Jokes/comments/3jwjrl/why_do_java_programmers_wear_glasses/,self.jokes,,because they can't C#,Why do Java programmers wear glasses?,165
post,3jwji7,2qh72,jokes,false,1441577754,https://old.reddit.com/r/Jokes/comments/3jwji7/if_i_got_a_dollar_everytime_someone_over_40_told/,self.jokes,,I'd have enough money to buy a house in the economy they ruined.,If I got a dollar everytime someone over 40 told me my generation sucks...,85
post,3jwjda,2qh72,jokes,false,1441577694,https://old.reddit.com/r/Jokes/comments/3jwjda/little_red_riding_hood/,self.jokes,,"Little red riding hood is walking in the forest when she hears a rustling in the bushes. She turns, and says “who’s there, oh who’s there?” Suddenly, the big bad wolf jumps up and runs off…

Later, little red is walking deeper in the woods and she hears a rustling in the bushes, so she turns and calls out again “who’s there, oh who’s there?”. Once again, the wolf jumps up and runs off into the bushes.

When Red riding hood is almost at her grandmothers, she hears another rustling in the bushes. Growing more anxious as to the wolf’s intentions, she calls out “I demand to know who is there!” 

The wolf jumps up and shouts back “can you give me a fucking minute I’ve been trying to have a shit for the last half hour!”",Little red riding hood,4
post,3jwism,2qh72,jokes,false,1441577423,https://old.reddit.com/r/Jokes/comments/3jwism/jack_off/,self.jokes,,"Two managers are going over their budget for the next year. After analyzing expenses and revenues, they come to the conclusion that they will have to lay off one of their two assistants, Jack or Jane.

They go back and forth but can't decide who to lay off. Finally, one manager decides that they should lay off the first person who gets up from their desk.

In the meantime, Jane is hard at work but suddenly gets a headache. She gets some aspirin from her desk drawer and gets up from her desk to get some water.


One of the managers gets up to break the bad news to Jane.

Manager: ""Jane, I need to talk to you. I've got a problem. I either need to lay you or Jack off...""

Jane:""Well, jack-off. I've got a headache.""
",Jack off...,1447
post,3jwhtr,2qh72,jokes,false,1441576950,https://old.reddit.com/r/Jokes/comments/3jwhtr/my_thesaurus_is_awful/,self.jokes,,"Not only that, it's also awful.",My thesaurus is awful.,120
post,3jwhix,2qh72,jokes,false,1441576793,https://old.reddit.com/r/Jokes/comments/3jwhix/memes/,self.jokes,,"http://imgur.com/qe7LBx5

there",memes,3
post,3jwgxz,2qh72,jokes,false,1441576496,https://old.reddit.com/r/Jokes/comments/3jwgxz/what_do_you_call_a_mexican_with_one_arm_shorter/,self.jokes,,not evennnn,What do you call a mexican with one arm shorter than the other?,0
post,3jwgjr,2qh72,jokes,false,1441576291,https://old.reddit.com/r/Jokes/comments/3jwgjr/did_you_hear_about_that_feminist_that_got_raped/,self.jokes,,[deleted],Did you hear about that feminist that got raped?,0
post,3jwg8b,2qh72,jokes,false,1441576130,https://old.reddit.com/r/Jokes/comments/3jwg8b/knock_knock/,self.jokes,,[deleted],Knock Knock!,0
post,3jwfwz,2qh72,jokes,false,1441575973,https://old.reddit.com/r/Jokes/comments/3jwfwz/whats_this_o/,self.jokes,,[deleted],What's this ? :-O,0
post,3jwfv1,2qh72,jokes,false,1441575947,https://old.reddit.com/r/Jokes/comments/3jwfv1/how_does_snoop_dogg_keep_his_shirts_so_white/,self.jokes,,BLE-YATCH!,How does Snoop Dogg keep his shirts so white?,0
post,3jwfn8,2qh72,jokes,false,1441575819,https://old.reddit.com/r/Jokes/comments/3jwfn8/knock_knock_whos_there_madame_madame_who/,self.jokes,,My damn foot's stuck in door!  Open up!,"Knock, knock. Who's there? Madame. Madame who?",0
post,3jwflw,2qh72,jokes,false,1441575802,https://old.reddit.com/r/Jokes/comments/3jwflw/whats_the_deal_with_arsenal_fans/,self.jokes,,"They're not British, they're not fans, we should call them plastics.",What's the deal with Arsenal fans?,0
post,3jwevy,2qh72,jokes,false,1441575477,https://old.reddit.com/r/Jokes/comments/3jwevy/a_chinese_man_walks_into_an_american_bank/,self.jokes,,"and sees the man in front of him exchanging some swiss francs into a good chunk of change. Remembering the leftover walk-around money from his vacation, he returns with roughly the same amount of francs the next week and asks the teller to exchange them.

Upon receiving a sum much smaller than anticipated, he demands to know why.

""Fluctuations.""

The teller says.

At this, the Chinese man turns red in the face and yells,

""Oh yeah? Well fruck you yankees too!""",A Chinese man walks into an American bank,2
post,3jwev3,2qh72,jokes,false,1441575467,https://old.reddit.com/r/Jokes/comments/3jwev3/never_fall_in_love_with_a_tennis_player/,self.jokes,,Love means nothing to them.,Never fall in love with a tennis player.,0
post,3jwe7v,2qh72,jokes,false,1441575159,https://old.reddit.com/r/Jokes/comments/3jwe7v/an_unassuming_man_takes_a_seat_at_a_stool_in_a_bar/,self.jokes,,"...The bartender walks up to him and asks what he'd like to drink. The man says he'd like a $25 martini. Before the bartender leaves the man stops him

""I bet you $50 that I remove my left eye and hold it in my hand."" 

The bartender agrees, and the man takes out his glass left eye and holds it in his hand.

""Let's do another,"" says the man. ""I bet you $250 that I can touch my right eye to my teeth.""

Once again, the bartender agrees, and so the man takes out his dentures and touches them to his right eye. The bartender is in disbelief.

""Last one,"" the man says. He walks across the bar, takes an empty glass from one of the tables, and puts it on the floor. He then walks back to the bartender. ""I bet you $10,000 that I can pee into that glass from here and make it without spilling a drop."" Well of course the bartender agrees. This man must surely be stupid for making a bet like that, he thinks.

The man unbuttons his trousers, grasps his penis in his hands and begins to pee. Immediately, he starts to flail around wildly, still going strong. Pee flies everywhere! It hits the bartender full force.

""Well, give me my thousand bucks,"" says the bartender, now giddy from happiness even though he was dripping in piss. He won $10,000 after all. So the man does without a bit of discontent. The bartender asks him why he isn't unhappy. 

""I'm a professional better,"" answers the man. ""You see that Chinese man over there? I bet him $1,000,000 that I'd pee on you and you'd be happy."" 
",An unassuming man takes a seat at a stool in a bar...,52
post,3jwe2j,2qh72,jokes,false,1441575091,https://old.reddit.com/r/Jokes/comments/3jwe2j/a_man_is_walking_on_the_beach/,self.jokes,,[deleted],A man is walking on the beach.,0
post,3jwdzv,2qh72,jokes,false,1441575053,https://old.reddit.com/r/Jokes/comments/3jwdzv/whats_the_speed_limit_of_sex/,self.jokes,,68... any faster and you'll eat it. ,What's the speed limit of sex?,1
post,3jwdi1,2qh72,jokes,false,1441574818,https://old.reddit.com/r/Jokes/comments/3jwdi1/why_do_women_wear_makeup_and_perfume/,self.jokes,,[deleted],Why do women wear makeup and perfume?,0
post,3jwdf5,2qh72,jokes,false,1441574784,https://old.reddit.com/r/Jokes/comments/3jwdf5/why_was_the_toilet_paper_in_east_germany_so/,self.jokes,,So every asshole would turn red.,Why was the toilet paper in East Germany so harshly?,4
post,3jwcd8,2qh72,jokes,false,1441574283,https://old.reddit.com/r/Jokes/comments/3jwcd8/three_oaps_are_sitting_in_a_retirement_home/,self.jokes,,[removed],Three OAP's are sitting in a retirement home discussing life,1
post,3jwcd4,2qh72,jokes,false,1441574280,https://old.reddit.com/r/Jokes/comments/3jwcd4/hey_guys_i_invented_a_new_word/,self.jokes,,Plagiarism.,"Hey guys, I invented a new word!",9
post,3jwbss,2qh72,jokes,false,1441574014,https://old.reddit.com/r/Jokes/comments/3jwbss/i_just_want_to_confirm_voip_on_nokia_lumia_521_is/,self.jokes,,[removed],I just want to confirm voip on Nokia Lumia 521 is terrible right?,1
post,3jwaqj,2qh72,jokes,false,1441573590,https://old.reddit.com/r/Jokes/comments/3jwaqj/why_did_the_police_assault_the_crowd/,self.jokes,,Because a-peppering them would make them sneeze!,Why did the police assault the crowd?,0
post,3jwak2,2qh72,jokes,false,1441573507,https://old.reddit.com/r/Jokes/comments/3jwak2/what_do_you_call_a_cheap_circumcision/,self.jokes,,A rip off!,What do you call a cheap circumcision?,44
post,3jwafu,2qh72,jokes,false,1441573452,https://old.reddit.com/r/Jokes/comments/3jwafu/that_thought_though/,self.jokes,,"A teacher is teaching a class and she sees that Johnny isn't paying attention, so she asks him, ""If there are three ducks sitting on a fence, and you shoot one, how many are left?"" Johnny says, ""None."" The teacher asks, ""Why?"" Johnny says, ""Because the shot scared them all off."" The teacher says, ""No, two, but I like how you're thinking."" Johnny asks the teacher, ""If you see three women walking out of an ice cream parlor, one is licking her ice cream, one is sucking her ice cream, and one is biting her ice cream, which one is married?"" The teacher says, ""The one sucking her ice cream."" Johnny says, ""No, the one with the wedding ring, but I like how you're thinking!",That thought though..,12
post,3jwaan,2qh72,jokes,false,1441573388,https://old.reddit.com/r/Jokes/comments/3jwaan/a_family_of_huntergatherers_sits_down_to_dinner/,self.jokes,,"The daughter, the youngest member of the family, complains, ""There's a hair in my soup!""

""Well,"" replies her father, the hunter of the household, ""technically, it's a rabbit.""",A family of hunter-gatherers sits down to dinner,4
post,3jw9tb,2qh72,jokes,false,1441573188,https://old.reddit.com/r/Jokes/comments/3jw9tb/mr_president_two_brazilian_soldiers_were_killed/,self.jokes,,[deleted],"""Mr. President, two Brazilian soldiers were killed yesterday in Iraq.""",0
post,3jw9oc,2qh72,jokes,false,1441573141,https://old.reddit.com/r/Jokes/comments/3jw9oc/how_many_american_rugby_fans_does_it_take_to/,self.jokes,,Both of them,How many american rugby fans does it take to change a lightbulb,719
post,3jw94y,2qh72,jokes,false,1441572877,https://old.reddit.com/r/Jokes/comments/3jw94y/why_is_the_ocean_salty/,self.jokes,,Because the land doesn't wave back,Why is the ocean salty?,50
post,3jw93b,2qh72,jokes,false,1441572851,https://old.reddit.com/r/Jokes/comments/3jw93b/a_dyslexic_man/,self.jokes,,A Dyslexic man walks into a bra.,A dyslexic man..,0
post,3jw917,2qh72,jokes,false,1441572821,https://old.reddit.com/r/Jokes/comments/3jw917/guests_are_like_fish/,self.jokes,,"After three days, you should probably get rid of them. ",Guests are like fish,1
post,3jw8s4,2qh72,jokes,false,1441572691,https://old.reddit.com/r/Jokes/comments/3jw8s4/i_heard_they_were_going_to_fine_bad_drivers_100/,self.jokes,,"That's bit sexist, isn't it? 
",I heard they were going to fine bad drivers $100 on the spot.,0
post,3jw8oz,2qh72,jokes,false,1441572645,https://old.reddit.com/r/Jokes/comments/3jw8oz/nsfw_i_asked_my_roommate_if_she_would_suck_my/,self.jokes,,The dirty cocksucker said no!,[NSFW] I asked my roommate if she would suck my cock after I cleaned it...,10
post,3jw850,2qh72,jokes,false,1441572347,https://old.reddit.com/r/Jokes/comments/3jw850/nsfw_whats_the_difference_in_your_mom_and_a/,self.jokes,,[deleted],[NSFW] What's the difference in your mom and a mosquito?,0
post,3jw7x3,2qh72,jokes,false,1441572236,https://old.reddit.com/r/Jokes/comments/3jw7x3/the_perfect_son/,self.jokes,,"A: I have the perfect son. 
B: Does he smoke? 
A: No, he doesn't. 
B: Does he drink whiskey? 
A: No, he doesn't. 
B: Does he ever come home late? 
A: No, he doesn't. 
B: I guess you really do have the perfect son. How old is he? 
A: He will be six months old next Wednesday.",The Perfect Son.,2
post,3jw6n7,2qh72,jokes,false,1441571586,https://old.reddit.com/r/Jokes/comments/3jw6n7/ring_hello_hi_honey_this_is_daddy_is_mommy_near/,self.jokes,,"""No Daddy. She's upstairs in the bedroom with Uncle Paul.""

After a brief pause, Daddy says, ""But honey, you don't have an Uncle Paul.""

""Oh yes I do, and he's upstairs in the room with Mommy, right now.""

Another brief pause... ""Uh, okay then, this is what I want you to do. Put the phone down on the table, run upstairs and knock on the bedroom door and shout to Mommy that Daddy's car just pulled into the driveway.""

""Okay Daddy, just a minute.""

A few minutes later the little girl comes back to the phone. ""I did it Daddy."" ""And what happened honey?"" he asked.

Well, Mommy got all scared, jumped out of bed with no clothes on and ran around screaming. She tripped over the rug, hit her head on the dresser and now she isn't moving at all!""

""Oh my God!!! What about your Uncle Paul?""

""He jumped out of the bed with no clothes on, too. He was all scared and he jumped out of the back window and into the swimming pool. But I guess he didn't know that you took out the water last week to clean it. He hit the bottom of the pool and I think he may be dead!""

There was a long pause, then Daddy says,

""Wait, swimming pool? Is this 486-5731?""","*RING* ""Hello?"", ""Hi honey. This is Daddy. Is Mommy near the phone?""",150
post,3jw6mo,2qh72,jokes,false,1441571578,https://old.reddit.com/r/Jokes/comments/3jw6mo/how_can_you_tell_if_balls_are_ticklish/,self.jokes,,[deleted],How can you tell if balls are ticklish?,10
post,3jw5hq,2qh72,jokes,false,1441571026,https://old.reddit.com/r/Jokes/comments/3jw5hq/the_picture_of_the_french_flag/,self.jokes,,http://i.imgur.com/cx13xBc.png,The picture of the french flag.,0
post,3jw57j,2qh72,jokes,false,1441570892,https://old.reddit.com/r/Jokes/comments/3jw57j/christiano_ronaldo_came_all_over_his_lovers_face/,self.jokes,,[deleted],Christiano Ronaldo came all over his lover's face...,0
post,3jw4xr,2qh72,jokes,false,1441570755,https://old.reddit.com/r/Jokes/comments/3jw4xr/a_lion_tamer_goes_to_see_a_psychologist/,self.jokes,,"
He explains: ""Doctor, I'm depressed. My emotional state is all over the place. I had a great idea for a new act - I was so excited and happy at first - the act seemed to be progressing so well - but then, it wouldn't seem to be working at all. It's been so full of up's and downs, I can barely keep track of myself"".

""What was the act?"" asked the doctor.

""Well, first - instead of using lions, the hook was that I instead used trained arctic bears.
First the 10 bears each grab a large cut-out letter, A to J, from a wall - and then arrange themselves alphabetically on stools on stage - much to the cheer of the audience. But each time exactly two and only two of the bears are always arranging themselves in the wrong order"".

The Doctor paused with thought - and then exclaimed:

""This sounds like a classic case of bi-polar disorder""",A lion tamer goes to see a psychologist...,0
post,3jw4jp,2qh72,jokes,false,1441570554,https://old.reddit.com/r/Jokes/comments/3jw4jp/so_travis_scott/,self.jokes,,[removed],So Travis Scott,1
post,3jw43d,2qh72,jokes,false,1441570331,https://old.reddit.com/r/Jokes/comments/3jw43d/two_muffins_are_in_an_oven/,self.jokes,,"The first muffin said: Wow, it's hot in here. 
The other muffin looked at the muffin: AHH! a talking muffin! 


-not mine, heard it from a friend when I was a kid and he apparently got it from tv",Two muffins are in an oven...,0
post,3jw37d,2qh72,jokes,false,1441569881,https://old.reddit.com/r/Jokes/comments/3jw37d/the_movie_iron_man_2/,self.jokes,,[deleted],The movie Iron Man 2...,0
post,3jw30g,2qh72,jokes,false,1441569775,https://old.reddit.com/r/Jokes/comments/3jw30g/a_new_energy_drink_called_f5_just_came_out_its/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jw30g/a_new_energy_drink_called_f5_just_came_out_its/,,"A new energy drink called F5 just came out, It's super refreshing!",15
post,3jw2j2,2qh72,jokes,false,1441569534,https://old.reddit.com/r/Jokes/comments/3jw2j2/the_normal_everyday_trent_richardson_would_have/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jw2j2/the_normal_everyday_trent_richardson_would_have/,,"The normal, everyday Trent Richardson would have cable...",0
post,3jw2ho,2qh72,jokes,false,1441569511,https://old.reddit.com/r/Jokes/comments/3jw2ho/thank_you_to_the_spanish_public_for/,self.jokes,,...rallying round and providing new headlines.,Thank you to the Spanish public for. ..,0
post,3jw1hb,2qh72,jokes,false,1441569041,https://old.reddit.com/r/Jokes/comments/3jw1hb/an_old_gay_man_dies/,self.jokes,,[deleted],An old gay man dies,2
post,3jw1ez,2qh72,jokes,false,1441569008,https://old.reddit.com/r/Jokes/comments/3jw1ez/عقارات_الشيخ_زايد/,self.jokes,,[removed],عقارات الشيخ زايد,1
post,3jw0w8,2qh72,jokes,false,1441568778,https://old.reddit.com/r/Jokes/comments/3jw0w8/late_one_night_a_man_is_driving_down_the_road/,self.jokes,,"Late one night a man is driving down the road, speeding quite a bit. A cop notices how fast he is going and pulls him over. The cop says to the man, ""Are you aware of how fast you were going?"" 

The man replies, ""Yes I am. I'm trying to escape a robbery I got involved in."" 

The cop gives him a skeptical look and says, ""Were you the one being robbed?"" 

The man casually replies, ""No, I committed the robbery."" 

The cop looks shocked that the man admitted this. ""So you're telling me you were speeding...AND committed a robbery?"" 

""Yes,"" the man calmly says. ""I have the loot in the back."" 

The cop begins to get angry. ""Sir, I'm afraid you have to come with me."" The cop reaches in the window to subdue the man. 

""Don't do that!"" the man yells fearfully. ""I'm scared you will find the gun in my glove compartment!"" The cop pulls his hand out. ""Wait here,"" he says. 

The cop calls for backup. Soon cops, cars, and helicopters are flooding the area. The man is cuffed quickly and taken towards a car. However, before he gets in, a cop walks up to him and says, while gesturing to the cop that pulled him over, ""Sir, this officer informed us that you had committed a robbery, had stolen loot in the trunk of your car, and had a loaded gun in your glove compartment. However, we found none of these things in your car."" 

The man replies, ""Yeah, and I bet that liar said I was speeding too!""","Late one night a man is driving down the road, speeding quite a bit...",10
post,3jvzis,2qh72,jokes,false,1441568009,https://old.reddit.com/r/Jokes/comments/3jvzis/an_irishman_a_scotsman_and_an_amnesiac_stumble/,self.jokes,,"The Irishman nearly escapes a speeding car, but the Scotsman isn't so lucky, and gets hit by the car and dies.","An Irishman, a Scotsman, and an amnesiac stumble drunkenly into the road.",3
post,3jvywl,2qh72,jokes,false,1441567743,https://old.reddit.com/r/Jokes/comments/3jvywl/how_do_you_starve_a_lazy_person/,self.jokes,,You put the welfare check in his work boots.,How do you starve a lazy person.,0
post,3jvyui,2qh72,jokes,false,1441567700,https://old.reddit.com/r/Jokes/comments/3jvyui/why_did_the_boy_drop_his_ice_cream/,self.jokes,,[deleted],Why did the boy drop his ice cream?,0
post,3jvyh4,2qh72,jokes,false,1441567512,https://old.reddit.com/r/Jokes/comments/3jvyh4/what_is_kurt_cobains_eye_color/,self.jokes,,"Blue. One blue to left, one blue to the right.",what is kurt cobain's eye color,0
post,3jvycn,2qh72,jokes,false,1441567448,https://old.reddit.com/r/Jokes/comments/3jvycn/what_do_you_call_the_place_where_a_bunch_of_nerds/,self.jokes,,[deleted],What do you call the place where a bunch of nerds hang out together because they have no place better to be?,0
post,3jvy87,2qh72,jokes,false,1441567391,https://old.reddit.com/r/Jokes/comments/3jvy87/a_pig_with_wings_walks_into_a_bar_stunned_the/,self.jokes,,"""You can't bring food in here from another restaurant! Even if you are a cop!""","A pig with wings walks into a bar. Stunned, the bartender says",200
post,3jvxht,2qh72,jokes,false,1441567066,https://old.reddit.com/r/Jokes/comments/3jvxht/whats_red_slime_and_crawls_up_your_leg/,self.jokes,,[deleted],"What's red, slime, and crawls up your leg?",0
post,3jvw8f,2qh72,jokes,false,1441566484,https://old.reddit.com/r/Jokes/comments/3jvw8f/epileptic_with_a_sword/,self.jokes,,"What do you get when an epileptic person fights an iceberg with a sword?

Seizure Salad",epileptic with a sword,0
post,3jvw40,2qh72,jokes,false,1441566431,https://old.reddit.com/r/Jokes/comments/3jvw40/what_do_you_get_when_you_break_a_babys_jaw/,self.jokes,,[deleted],What do you get when you break a baby's jaw?,0
post,3jvvy6,2qh72,jokes,false,1441566354,https://old.reddit.com/r/Jokes/comments/3jvvy6/how_do_chinese_officials_get_elected_to_office/,self.jokes,,[deleted],How do Chinese officials get elected to office?,0
post,3jvvs1,2qh72,jokes,false,1441566269,https://old.reddit.com/r/Jokes/comments/3jvvs1/what_arent_drunken_noodles/,self.jokes,,[deleted],What aren't drunken noodles?,0
post,3jvvlt,2qh72,jokes,false,1441566185,https://old.reddit.com/r/Jokes/comments/3jvvlt/now_that_i_downloaded_true_caller_i_hope_i_find/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jvvlt/now_that_i_downloaded_true_caller_i_hope_i_find/,,"Now that I downloaded True Caller, I hope I find my true calling.",0
post,3jvv8z,2qh72,jokes,false,1441566021,https://old.reddit.com/r/Jokes/comments/3jvv8z/whats_chinese_and_climbs_the_empire_state_building/,self.jokes,,Ping Pong,What's Chinese and climbs the Empire State Building?,1
post,3jvup0,2qh72,jokes,false,1441565770,https://old.reddit.com/r/Jokes/comments/3jvup0/why_was_the_energizer_bunny_arrested/,self.jokes,,He was charged with battery. XD,Why was the Energizer Bunny arrested?,1
post,3jvuly,2qh72,jokes,false,1441565736,https://old.reddit.com/r/Jokes/comments/3jvuly/three_professors_go_to_the_nudist_beach/,self.jokes,,"They start reading their newspapers, when suddenly Miss Ridgewell approaches them from the Chemistry Department. The alarmed professors react immediately. Two of them hide their manhood with their newspapers, the third, however, hides his face. They politely salute the lady, who simply passes by to join her friends.

When she's far gone, one of them asks the third professor, ""Why did you hide your face?""

To which the third professor replies, ""I don't know about you guys, but people usually recognise my face...""",Three professors go to the nudist beach,36
post,3jvu4l,2qh72,jokes,false,1441565526,https://old.reddit.com/r/Jokes/comments/3jvu4l/two_fish_in_a_tank/,self.jokes,,"Fish 1: uh, Greg?


Fish 2: what


Fish 1: how do we drive this thing",Two fish in a tank,40
post,3jvtmw,2qh72,jokes,false,1441565301,https://old.reddit.com/r/Jokes/comments/3jvtmw/jesus_take_the_wheel/,self.jokes,,"Carlos you take the stereo
I'll take lookout ",Jesus take the wheel,464
post,3jvsyh,2qh72,jokes,false,1441565003,https://old.reddit.com/r/Jokes/comments/3jvsyh/my_friend_is_like_a_jew_during_wwii/,self.jokes,,In the closet.,My friend is like a Jew during WWII,1
post,3jvsv2,2qh72,jokes,false,1441564955,https://old.reddit.com/r/Jokes/comments/3jvsv2/a_doctor_on_his_morning_walk_noticed_an_old_lady/,self.jokes,,"A doctor on his morning walk noticed an old lady sitting on her front step smoking a cigar 



So he walked up to her and said, ""I couldn't help but notice how happy you look! What is your secret?"" 




""I smoke ten cigars a day,"" she said. '""Before I go to bed, I smoke a nice big joint. Apart from that, I drink a whole bottle of Jack Daniels every week, and eat only junk food. On weekends, I pop pills, get laid, and don't exercise at all.""



'""That is absolutely amazing! How old are you?""



""Thirty-four,"" she replied. ",A doctor on his morning walk noticed an old lady sitting on her front step smoking a cigar,39
post,3jvsu6,2qh72,jokes,false,1441564944,https://old.reddit.com/r/Jokes/comments/3jvsu6/one_day_in_the_great_forest_a_magical_frog_was/,self.jokes,,[deleted],"One day in the great forest, a magical frog was walking down to a water hole.",6
post,3jvsn6,2qh72,jokes,false,1441564858,https://old.reddit.com/r/Jokes/comments/3jvsn6/i_eat_more_pussy_than_cervical_cancer_nsfw/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jvsn6/i_eat_more_pussy_than_cervical_cancer_nsfw/,,I eat more pussy than cervical cancer. [NSFW],0
post,3jvr9c,2qh72,jokes,false,1441564250,https://old.reddit.com/r/Jokes/comments/3jvr9c/whats_common_between_a_lawyer_and_an_eccentric/,self.jokes,,Both have a very expensive retainer.,What's common between a lawyer and an eccentric billionaire with bad teeth?,2
post,3jvr6g,2qh72,jokes,false,1441564216,https://old.reddit.com/r/Jokes/comments/3jvr6g/nsfw_i_eat_more_pussy_than_cervical_cancer/,self.jokes,,[deleted],NSFW I eat more pussy than cervical cancer.,1
post,3jvqv6,2qh72,jokes,false,1441564008,https://old.reddit.com/r/Jokes/comments/3jvqv6/one_of_my_freind_like_this_joke/,self.jokes,,"hey bro,Today a  man knocked on my door and asked for a small donation towards the local swimming pool.

cool,so did you help him bro?

yes bro,i gave him a glass of water.
",one of my freind like this joke.,1
post,3jvqse,2qh72,jokes,false,1441563973,https://old.reddit.com/r/Jokes/comments/3jvqse/what_do_you_get_if_you_mix_a_joke_with_a/,self.jokes,,[deleted],What do you get if you mix a joke with a rhetorical question?,1
post,3jvqsb,2qh72,jokes,false,1441563973,https://old.reddit.com/r/Jokes/comments/3jvqsb/why_is_it_so_hard_for_an_eighty_year_old_woman_to/,self.jokes,,Have you ever tried pulling apart a grilled cheese?!,Why is it so hard for an eighty year old woman to pee in the morning?,0
post,3jvphu,2qh72,jokes,false,1441563389,https://old.reddit.com/r/Jokes/comments/3jvphu/fishing/,self.jokes,,Give a kid a fish he can eat for a day. Teach a kid to fish he can eat for life. Give him a fishing rod he can find his dad at the bottom of a lake in Syria,Fishing,0
post,3jvotb,2qh72,jokes,false,1441563084,https://old.reddit.com/r/Jokes/comments/3jvotb/im_friends_with_25_letters_of_the_alphabet/,self.jokes,,"I don´t know y



DDD",i´m friends with 25 letters of the alphabet,2
post,3jvnz4,2qh72,jokes,false,1441562710,https://old.reddit.com/r/Jokes/comments/3jvnz4/my_favorite_joke_to_play_on_people_with_stretched/,self.jokes,,[deleted],My favorite joke to play on people with stretched ear holes/plugs/GUAGES... works like a charm! :),0
post,3jvnbg,2qh72,jokes,false,1441562400,https://old.reddit.com/r/Jokes/comments/3jvnbg/a_stick_figure_walks_into_a_bar_and_takes_five/,self.jokes,,He's dead.,"A stick figure walks into a bar, and takes five shots.",0
post,3jvm22,2qh72,jokes,false,1441561803,https://old.reddit.com/r/Jokes/comments/3jvm22/how_do_nazis_measure_the_intensity_of_earthquakes/,self.jokes,,[deleted],How do Nazis measure the intensity of earthquakes?,1
post,3jvm1d,2qh72,jokes,false,1441561793,https://old.reddit.com/r/Jokes/comments/3jvm1d/why_was_the_smurfs_hat_blue/,self.jokes,,Cus it was sad.,Why was the smurf's hat blue?,0
post,3jvl01,2qh72,jokes,false,1441561293,https://old.reddit.com/r/Jokes/comments/3jvl01/what_is_the_politically_correct_term_for_middle/,self.jokes,,[deleted],What is the Politically Correct term for Middle Easterners in the U.S.?,0
post,3jvkpl,2qh72,jokes,false,1441561152,https://old.reddit.com/r/Jokes/comments/3jvkpl/i_opened_the_window/,self.jokes,,And influenza.,I opened the window...,3
post,3jvke1,2qh72,jokes,false,1441561004,https://old.reddit.com/r/Jokes/comments/3jvke1/nymphomaniac_convention/,self.jokes,,"I have no idea if this has been posted here before, so I apologize if it's a repost, otherwise enjoy.

A man is boarding plane to Vegas when a very attractive young woman takes the seat next to him. They start talking about various things, and he asks why  she's going to Las Vegas, and is very surprised to hear that she intends to give a lecture at the annual Nymphomaniac Convention.

After he inquires what she plans to lecture about, she tells him she is going to attempt to dispel a few sexual myths and attempt to give some much needed insight to the people of America. Utterly intrigued, he listens as she tells him that it is, in fact, not African Americans who are the most well endowed, but Native Americans. Though it is usually believed that the French are among the most skilled lovers, the Jewish actually tend to be even better. The least expected thing she said though was that the typical southern redneck had the best stamina of any other  typical profile or stereotype out there.

As the man is sitting there just taking it all in, the woman realizes she's been going on and on about her interests and doesn't even know his name yet, so she asks him, to which he replies ""My name? Tonto, Tonto Goldstein, but my friends call me Bubba.""",Nymphomaniac Convention,0
post,3jvjuy,2qh72,jokes,false,1441560760,https://old.reddit.com/r/Jokes/comments/3jvjuy/why_is_lemon_juice_made_with_artificial_flavor/,self.jokes,,[deleted],"Why is lemon juice made with artificial flavor, and dishwashing liquid made with real lemons . Why is the alphabet in that order?",0
post,3jvjjg,2qh72,jokes,false,1441560586,https://old.reddit.com/r/Jokes/comments/3jvjjg/on_a_scale_of_110_how_funny_is_reddit/,self.jokes,,Probably banana ,"on a scale of 1-10, how funny is reddit?",1
post,3jviym,2qh72,jokes,false,1441560320,https://old.reddit.com/r/Jokes/comments/3jviym/a_man_taking_on_a_late_night_walk_when_he_hears_a/,self.jokes,,"As he approaches he realizes he's hearing chanting. He approaches the building and hears ""sixty-seven! Sixty-seven! Sixty-seven!"" He gets closer to investigate but the fence is too high to see over, though he does spot a small hole in the wood. He leans over to peep in and as soon as he does a finger pokes him in the eye, and he hears the man on the other end shout ""sixty-eight!""",A man taking on a late night walk when he hears a strange sound coming from an old mental hospital down the road.,8
post,3jvis7,2qh72,jokes,false,1441560234,https://old.reddit.com/r/Jokes/comments/3jvis7/how_come_mr_and_mrs_claus_dont_have_any_kids/,self.jokes,,Because Santa only cums once a year and its down the chimney!,How come Mr. and Mrs. Claus don't have any kids?,23
post,3jvior,2qh72,jokes,false,1441560189,https://old.reddit.com/r/Jokes/comments/3jvior/a_little_boy_aged_7_asks_dad_daddy_what_is_sex/,self.jokes,,"Shocked by his son's question , dad felt that he shouldn't lie to his son . Dad began ,"" son when a man and woman ..."" After a detailed explanation dad finished. Then his son replied ,""Daddy mom said that breakfast will be ready in 60 sex ( secs ) .","A little boy , aged 7 asks dad , ""daddy what is sex "" ?",1
post,3jvinn,2qh72,jokes,false,1441560173,https://old.reddit.com/r/Jokes/comments/3jvinn/why_did_the_baker_have_sticky_hands/,self.jokes,,Because he kneaded a poo.,Why did the baker have sticky hands?,0
post,3jvihq,2qh72,jokes,false,1441560095,https://old.reddit.com/r/Jokes/comments/3jvihq/a_philosopher_walks_into_a_bank_and_exclaims/,self.jokes,,[deleted],A philosopher walks into a bank and exclaims...,0
post,3jvig2,2qh72,jokes,false,1441560076,https://old.reddit.com/r/Jokes/comments/3jvig2/gave_my_wife_a_coffee_enema/,self.jokes,,"Gave my wife a coffee enema. She grimaced. I asked, ""too hot""? ""No"", she replied, ""too sweet"".",Gave my wife a coffee enema,0
post,3jvi75,2qh72,jokes,false,1441559961,https://old.reddit.com/r/Jokes/comments/3jvi75/what_do_9_out_of_10_people_enjoy/,self.jokes,,Gang rape.,What do 9 out of 10 people enjoy?,1
post,3jvha0,2qh72,jokes,false,1441559508,https://old.reddit.com/r/Jokes/comments/3jvha0/whats_a_single_mothers_favorite_dessert/,self.jokes,,creampie ,What's a single mother's favorite dessert?,2
post,3jvgm9,2qh72,jokes,false,1441559199,https://old.reddit.com/r/Jokes/comments/3jvgm9/what_did_david_say_when_the_tourist_tried_to/,self.jokes,,Don't touch my marbles.,What did David say when the tourist tried to touch him?,0
post,3jvglx,2qh72,jokes,false,1441559195,https://old.reddit.com/r/Jokes/comments/3jvglx/the_canadian_army/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jvglx/the_canadian_army/,,The Canadian Army,0
post,3jvggc,2qh72,jokes,false,1441559114,https://old.reddit.com/r/Jokes/comments/3jvggc/cooking_hack/,self.jokes,,[deleted],COOKING HACK,2
post,3jvgej,2qh72,jokes,false,1441559091,https://old.reddit.com/r/Jokes/comments/3jvgej/why_cant_your_penis_be_12_inches/,self.jokes,,Because then it'd be a foot,Why can't your penis be 12 inches?,9
post,3jvfog,2qh72,jokes,false,1441558736,https://old.reddit.com/r/Jokes/comments/3jvfog/wanna_hear_a_good_pickup_line/,self.jokes,,[deleted],Wanna hear a good pickup line?,0
post,3jvf4d,2qh72,jokes,false,1441558473,https://old.reddit.com/r/Jokes/comments/3jvf4d/how_does_a_train_driver_operate_a_train_while/,self.jokes,,"He goes chew chew chew...


creds to my 5yo brother",How does a train driver operate a train while eating gum?,14
post,3jveld,2qh72,jokes,false,1441558234,https://old.reddit.com/r/Jokes/comments/3jveld/does_anyone_know_what_subreddit_your_mamma_jokes/,self.jokes,,Jk. ,"Does anyone know what subreddit ""your mamma"" jokes are in?",0
post,3jvdfg,2qh72,jokes,false,1441557679,https://old.reddit.com/r/Jokes/comments/3jvdfg/why_should_you_never_bet_on_germany_at_the/,self.jokes,,They have the worst track record for finishing a race.,Why should you never bet on Germany at the Olympics?,0
post,3jvctc,2qh72,jokes,false,1441557393,https://old.reddit.com/r/Jokes/comments/3jvctc/little_johnny/,self.jokes,,"Little Johnny is in the first grade and learning the letters of the alphabet.  His teacher is calling on students to tell her a word that starts with each letter.  When she asks for a word that starts with A, immediately Johnny raises his hand.  Now, the teacher knows he is going to say something dirty like asshole so she won't call on him.  Same thing for the letter B.  Johnny raises his hand but the teacher is afraid he'll say bitch or boobs.  This goes on for almost the entire alphabet until they get to the letter ""R"".  The teacher can't think of anything dirty so she goes ahead and calls on Johnny.  He then says, ""Rabbit"".  The teacher starts to tell him that this is very nice answer, but Johnny cuts her off by saying ""WITH A COCK THIS FUCKING BIG!"" ",Little Johnny...,3
post,3jvcpy,2qh72,jokes,false,1441557346,https://old.reddit.com/r/Jokes/comments/3jvcpy/a_jewish_boy_asks_his_father/,self.jokes,,"A Jewish boy asks his Father, ""Dad, can i have 50 pence please?

His Father replies, ""40 pence! What do you want 30 pence for?""",A Jewish boy asks his Father...,10
post,3jvc64,2qh72,jokes,false,1441557067,https://old.reddit.com/r/Jokes/comments/3jvc64/is_it_wrong_to_hate_a_certain_race/,self.jokes,,Because I despise the 200 meter sprint.,is it wrong to hate a certain race?,1
post,3jvbxv,2qh72,jokes,false,1441556952,https://old.reddit.com/r/Jokes/comments/3jvbxv/babe_some_guy_told_me_today_that_if_i_have_sex/,self.jokes,,... he'll give me these earrings. What a jerk!,"Babe, some guy told me today that if I have sex with him...",0
post,3jvbt0,2qh72,jokes,false,1441556885,https://old.reddit.com/r/Jokes/comments/3jvbt0/why_does_youtube_have_a_stable_ph/,self.jokes,,'Cause it buffers a lot.,Why does YouTube have a stable pH??,1
post,3jvbma,2qh72,jokes,false,1441556792,https://old.reddit.com/r/Jokes/comments/3jvbma/if_you_have_dad_issues/,self.jokes,,[deleted],If you have dad issues...,0
post,3jvbfa,2qh72,jokes,false,1441556690,https://old.reddit.com/r/Jokes/comments/3jvbfa/how_do_you_find_will_smith_in_a_snow_storm/,self.jokes,,Follow the fresh prints ,How do you find will smith in a snow storm?,21
post,3jvbam,2qh72,jokes,false,1441556636,https://old.reddit.com/r/Jokes/comments/3jvbam/a_woman_brings_her_elderly_husband_to_the_doctor/,self.jokes,,"A woman brings her elderly husband to the doctor for his annual check-up.  After the examination, the doctor pulls the woman aside.

""Your husband is in good physical shape,"" he says, ""But I'm concerned about his mental health.  He told me that when he gets up to go to the bathroom at night, God turns on the light for him.""

""Oh, damn!"" the wife replies, ""He's pissing in the refrigerator again.""",A woman brings her elderly husband to the doctor for his annual check-up.,102
post,3jvb6y,2qh72,jokes,false,1441556586,https://old.reddit.com/r/Jokes/comments/3jvb6y/i_am_the_walruskukukajoo/,self.jokes,,"Q: Why did the Walrus go to the Tupperware Party?

A: he was looking for a Tight-Seal",I am the Walrus....ku-ku-ka-joo,1
post,3jvb4o,2qh72,jokes,false,1441556555,https://old.reddit.com/r/Jokes/comments/3jvb4o/where_does_monty_python_buy_his_water/,self.jokes,,"From the knights Da-sa(y)-NI! 


This joke is best delivered verbally.

",Where does monty python buy his water?,0
post,3jvaxw,2qh72,jokes,false,1441556463,https://old.reddit.com/r/Jokes/comments/3jvaxw/what_does_time_do_when_its_still_hungry/,self.jokes,,[deleted],What does time do when it's still hungry?,3
post,3jvany,2qh72,jokes,false,1441556333,https://old.reddit.com/r/Jokes/comments/3jvany/the_number/,self.jokes,,"One day,i saw a girl whose Facebook name is 70.Because of curiosity I added her.Until i have done with her and her name changed to 71, i know what her means.",The number,0
post,3jva1k,2qh72,jokes,false,1441556026,https://old.reddit.com/r/Jokes/comments/3jva1k/dad_joke_what_do_you_get_when_you_combine_a/,self.jokes,,[removed],Dad Joke: What do you get when you combine a computer with an elephant?,1
post,3jv8t9,2qh72,jokes,false,1441555433,https://old.reddit.com/r/Jokes/comments/3jv8t9/my_roommate_just_called_my_clothes_gay/,self.jokes,,Have a little respect man! They just came out of the closet,My roommate just called my clothes gay..,360
post,3jv8oc,2qh72,jokes,false,1441555373,https://old.reddit.com/r/Jokes/comments/3jv8oc/why_do_jews_play_football/,self.jokes,,So they can get the Quarterback!,Why Do Jews Play Football?,0
post,3jv8fz,2qh72,jokes,false,1441555248,https://old.reddit.com/r/Jokes/comments/3jv8fz/what_happened_to_the_number_10/,self.jokes,,It got stuck in 9/11,What happened to the number 10?,1
post,3jv7am,2qh72,jokes,false,1441554708,https://old.reddit.com/r/Jokes/comments/3jv7am/whats_a_pirates_favorite_letter/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jv7am/whats_a_pirates_favorite_letter/,,What's a pirate's favorite letter?,1
post,3jv6v4,2qh72,jokes,false,1441554499,https://old.reddit.com/r/Jokes/comments/3jv6v4/i_ran_into_my_x_the_other_day/,self.jokes,, Now I have to get my bicycle repaired.,I ran into my X the other day.,1
post,3jv62u,2qh72,jokes,false,1441554111,https://old.reddit.com/r/Jokes/comments/3jv62u/during_last_nights_couples_massage_my_female/,self.jokes,," both massage therapist are blown away. All I can think is my wife  &amp;  boss ride my back 24/7. This is easy.

 #RealLife  
PS: My helicopter boss and wife share the same name. 
#MarriedLife4Lyfe","During last nights couples massage, my female masseuse mounts my back with full weight on her knees and......",0
post,3jv5uu,2qh72,jokes,false,1441553989,https://old.reddit.com/r/Jokes/comments/3jv5uu/whats_the_difference_between_911_and_a_cow/,self.jokes,,[deleted],What's the difference between 9/11 and a cow?,0
post,3jv5lg,2qh72,jokes,false,1441553848,https://old.reddit.com/r/Jokes/comments/3jv5lg/why_do_all_chinese_planes_have_treasure_chests_on/,self.jokes,,Because they are flown by Pirots.  (Pirates),Why do all Chinese planes have treasure chests on board?,0
post,3jv5im,2qh72,jokes,false,1441553803,https://old.reddit.com/r/Jokes/comments/3jv5im/what_does_a_mafioso_and_rick_astley_have_in_common/,self.jokes,,They're never going to give you up. ,What does a Mafioso and Rick Astley have in common?,0
post,3jv4rb,2qh72,jokes,false,1441553403,https://old.reddit.com/r/Jokes/comments/3jv4rb/why_are_pills_white/,self.jokes,,[deleted],Why are pills white?,0
post,3jv4kp,2qh72,jokes,false,1441553295,https://old.reddit.com/r/Jokes/comments/3jv4kp/a_family_walks_into_a_hotel/,self.jokes,,"A family walks into a hotel and the father goes to the front desk and says ""I hope the porn is disabled."" The guy at the desk replies ""it's just regular porn, you sick fuck.""  ",A family walks into a hotel...,61
post,3jv4j4,2qh72,jokes,false,1441553277,https://old.reddit.com/r/Jokes/comments/3jv4j4/my_friend_said_when_my_mum_was_pregnant_with_me/,self.jokes,,[deleted],"My friend said, ""When my mum was pregnant with me she was very sick""",0
post,3jv46y,2qh72,jokes,false,1441553093,https://old.reddit.com/r/Jokes/comments/3jv46y/how_many_statisticians_does_it_take_to_screw_a/,self.jokes,,[deleted],How many statisticians does it take to screw a light bulb?,0
post,3jv43m,2qh72,jokes,false,1441553049,https://old.reddit.com/r/Jokes/comments/3jv43m/pulled_up_next_to_a_guy_with_a_new_england/,self.jokes,,[deleted],Pulled up next to a guy with a New England Patriots bumper sticker...,0
post,3jv3lp,2qh72,jokes,false,1441552818,https://old.reddit.com/r/Jokes/comments/3jv3lp/i_could_tell_you_that_sodium_hydroxide_is_a/,self.jokes,,But then that would be a lye.,I could tell you that sodium hydroxide is a liquid out of solution.,43
post,3jv3ah,2qh72,jokes,false,1441552643,https://old.reddit.com/r/Jokes/comments/3jv3ah/my_dentist_took_a_look_in_my_mouth_and_said_your/,self.jokes,,"I do, I said, I floss on Christmas and Easter.","My dentist took a look in my mouth and said, ""Your gums look awful. I told you to floss religiously.""",26
post,3jv359,2qh72,jokes,false,1441552576,https://old.reddit.com/r/Jokes/comments/3jv359/a_boy_tells_his_father_hes_lost_his_virginity/,self.jokes,,[deleted],A boy tells his father he's lost his virginity,0
post,3jv2xl,2qh72,jokes,false,1441552471,https://old.reddit.com/r/Jokes/comments/3jv2xl/what_is_the_difference_between_your_gullibility/,self.jokes,,[deleted],What is the difference between your gullibility and the punchline of this joke?,0
post,3jv299,2qh72,jokes,false,1441552128,https://old.reddit.com/r/Jokes/comments/3jv299/john_get_angry/,self.jokes,,"So John is standing on a bus stop waiting for bus.
In meantime, a woman with kid comes to wait for bus aswell.
As any other kid, this kid gets restless and ask mom: 
-why is bus not here yet moma
Mom replies:
- they are washing it honey.
After few minutes kid asks again:
-mommy, why is bus not here yet?
-They are fixing the engine hon.
Minutes later kid asks again:
-why is bus still not here mom?
-They are doing a paint job sweaty.
Hearing that John bursts in rage :
- Do THEY seriously thik that now is the best time to start painting their bus??????",John get angry,0
post,3jv1f5,2qh72,jokes,false,1441551704,https://old.reddit.com/r/Jokes/comments/3jv1f5/what_do_you_call_a_stupid_robot/,self.jokes,,[deleted],What do you call a stupid robot?,1
post,3jv16z,2qh72,jokes,false,1441551595,https://old.reddit.com/r/Jokes/comments/3jv16z/in_russia_if_youre_blue_and_you_dont_where_to_go/,self.jokes,,Putin on the Ritz,"In Russia, if you're blue, and you don't where to go to, why don't you go where fashion sits:",0
post,3juztf,2qh72,jokes,false,1441550862,https://old.reddit.com/r/Jokes/comments/3juztf/man_arrives_home_at_7_am_with_a_heavy_stench_of/,self.jokes,,"Wife: You bastard! I hope you have a damn good reason for coming home at 7 in the morning. 

Husband: Of course I do.

Wife: Do tell!

Husband: Breakfast.","Man arrives home at 7 a.m, with a heavy stench of whisky.",1304
post,3juzs5,2qh72,jokes,false,1441550843,https://old.reddit.com/r/Jokes/comments/3juzs5/women_are_like_farts/,self.jokes,,[deleted],Women are like farts...,0
post,3juzpk,2qh72,jokes,false,1441550804,https://old.reddit.com/r/Jokes/comments/3juzpk/my_grandfather_was_extremely_proud_of_his/,self.jokes,,[deleted],"My grandfather was extremely proud of his completely British heritage, but then he found out his grandmother actually came from Transylvania.",3
post,3juytm,2qh72,jokes,false,1441550314,https://old.reddit.com/r/Jokes/comments/3juytm/what_did_the_buddhist_say_to_the_hot_dog_vendor/,self.jokes,,[removed],What did the Buddhist say to the hot dog vendor?,0
post,3juyem,2qh72,jokes,false,1441550074,https://old.reddit.com/r/Jokes/comments/3juyem/i_went_shopping_with_my_wife_the_other_day_and/,self.jokes,,[deleted],I went shopping with my wife the other day and after entering the store she called me fat and lazy,4
post,3juy9x,2qh72,jokes,false,1441549987,https://old.reddit.com/r/Jokes/comments/3juy9x/an_elderly_woman_is_discussing_genderroles_with/,self.jokes,,[deleted],An elderly woman is discussing gender-roles with her granddaughter.,0
post,3juy5s,2qh72,jokes,false,1441549911,https://old.reddit.com/r/Jokes/comments/3juy5s/hey/,self.jokes,,Click this link. ,Hey,0
post,3juxjm,2qh72,jokes,false,1441549554,https://old.reddit.com/r/Jokes/comments/3juxjm/watch_and_enjoy_vid/,self.jokes,,[removed],Watch and enjoy (vid),1
post,3jux9s,2qh72,jokes,false,1441549422,https://old.reddit.com/r/Jokes/comments/3jux9s/two_midgets_decide_to_get_hookers/,self.jokes,,"They went to a motel with their ladies and get two rooms.  The first midget is really embarrassed because he cannot get an erection.  His confidence was hurt even more when he heard his friend in the room saying ""1, 2, 3, push!"" Over and over again.

The next morning he was talking to his friend over breakfast. He said ""That was the most embarrassing thing ever.  I couldn't get a hard on""
His friend responds ""You think that is embarrassing, I couldn't get on the bed.""

Edit:spelling ",Two midgets decide to get hookers...,46
post,3jux7i,2qh72,jokes,false,1441549374,https://old.reddit.com/r/Jokes/comments/3jux7i/a_soldier_wakes_up_one_morning/,self.jokes,,"A soldier wakes up one morning and goes down to breakfast. He has tousled hair and deep, dark bags under his eyes. 

""How did you sleep, honey?"" his mom asks. 

""Like Iraq,"" he answers. 

""That's great, sweetie,"" she says without looking up. ",A soldier wakes up one morning...,2
post,3jux3i,2qh72,jokes,false,1441549306,https://old.reddit.com/r/Jokes/comments/3jux3i/i_decided_not_to_go_on_that_date_with_the_bank/,self.jokes,,No interest,I decided not to go on that date with the bank teller,2
post,3jux0l,2qh72,jokes,false,1441549254,https://old.reddit.com/r/Jokes/comments/3jux0l/a_green_man_is_having_a_shower/,self.jokes,,"...a woman knocks on the door, the man wraps a towel around himself and answers it. They start to have a conversation then the mans towel falls down. The woman screams, runs off and is hit by a car. Moral of the story: never run when the green man's flashing. ",A green man is having a shower...,1
post,3juwm8,2qh72,jokes,false,1441549000,https://old.reddit.com/r/Jokes/comments/3juwm8/mickey_mouse_and_minnie_mouse_are_getting_a/,self.jokes,,"Mickey Mouse and Minnie Mouse are getting a divorce. The judge says to Mickey, ""Mr. Mouse, for the last time, I'm trying to explain to you that you can't divorce Minnie because she's stupid."" Mickey says, ""Your honor, for the last time, I don't want to divorce Minnie because she's stupid, I want to divorce her because she's fucking Goofy.""",Mickey Mouse and Minnie Mouse are getting a divorce,3
post,3juwi7,2qh72,jokes,false,1441548936,https://old.reddit.com/r/Jokes/comments/3juwi7/why_was_6_afraid_of_7/,self.jokes,,Because 7 was a registered 6 offender.,Why was 6 afraid of 7?,69
post,3juwah,2qh72,jokes,false,1441548807,https://old.reddit.com/r/Jokes/comments/3juwah/what_do_you_call_a_wellendowed_member_of_hitlers/,self.jokes,,Hungaryan.,What do you call a well-endowed member of Hitler's master race?,9
post,3juw2d,2qh72,jokes,false,1441548674,https://old.reddit.com/r/Jokes/comments/3juw2d/despite_the_large_variations_in_ambient/,self.jokes,,By definition.,"Despite the large variations in ambient temperature, how do warm blooded animals stay warm?",0
post,3juvua,2qh72,jokes,false,1441548541,https://old.reddit.com/r/Jokes/comments/3juvua/what_do_you_call_a_wellendowed_member_of_hitlers/,self.jokes,,[deleted],What do you call a well-endowed member of Hitler's master race?,2
post,3juvj0,2qh72,jokes,false,1441548350,https://old.reddit.com/r/Jokes/comments/3juvj0/did_you_hear_about_the_constipated_chancellor/,self.jokes,,"He couldn't budge it :P

",Did you hear about the constipated chancellor?,7
post,3juvhy,2qh72,jokes,false,1441548336,https://old.reddit.com/r/Jokes/comments/3juvhy/the_kindness_of_strangers/,self.jokes,,"An old lady on a bus offers the driver some peanuts. The driver, being polite, accepts and munches them.

Every 5 minutes she gives him a handful more peanuts.

Driver : Why don't you eat them yourself ?

Old lady : I can't chew them. Look, I have no teeth.

Driver : Then why do you buy them ?

Old lady : Oh, I just love the chocolates around them.",The kindness of strangers,261
post,3juv9a,2qh72,jokes,false,1441548194,https://old.reddit.com/r/Jokes/comments/3juv9a/my_poem/,self.jokes,,"I dig...
You dig...
We dig...
He digs...
She digs...
They dig...
Now it's not a very beautiful poem, but it's quite deep",My poem,165
post,3juv11,2qh72,jokes,false,1441548065,https://old.reddit.com/r/Jokes/comments/3juv11/a_guy_and_a_girl_have_a_conversation_during_sex/,self.jokes,,"The guy says, ""So when's your birthday?""

The girl replies ""July 23rd.""

The guy says ""No way, me too!""

The girl gets excited and asks, ""No way, are you fucking with me?""

The guy looks down at his penis inserted in the girl's vagina and says, ""Well, technically, yes.""",A guy and a girl have a conversation during sex.,0
post,3jutyo,2qh72,jokes,false,1441547432,https://old.reddit.com/r/Jokes/comments/3jutyo/family_cat_had_severe_blood_loss/,self.jokes,,"The family cat had just suffered a horrific accident and had severe blood loss.  We brought the cat to the vet, who said that the only way to save our pet was to donate blood.  Luckily, we read over the medical papers and it was type AB so anyone could donate blood; I volunteered.  The doctor performed the procedure, but alas the cat died.  Turned out, it was a typo.",Family cat had severe blood loss...,1
post,3jutvg,2qh72,jokes,false,1441547376,https://old.reddit.com/r/Jokes/comments/3jutvg/kim_davis/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jutvg/kim_davis/,,Kim Davis,0
post,3jutgt,2qh72,jokes,false,1441547107,https://old.reddit.com/r/Jokes/comments/3jutgt/a_family_walks_into_a_talent_agency/,self.jokes,,[removed],A family walks into a talent agency,0
post,3jut47,2qh72,jokes,false,1441546880,https://old.reddit.com/r/Jokes/comments/3jut47/why_do_skeletons_not_go_to_the_disco/,self.jokes,,Because they got no body to dance with!,Why do skeletons not go to the disco?,5
post,3jusgi,2qh72,jokes,false,1441546447,https://old.reddit.com/r/Jokes/comments/3jusgi/a_family_walks_into_a_talent_agency/,self.jokes,,[removed],A family walks into a talent agency,1
post,3jurni,2qh72,jokes,false,1441545923,https://old.reddit.com/r/Jokes/comments/3jurni/which_is_worse_ignorance_or_apathy/,self.jokes,,I don't know and I don't care.,Which is worse: ignorance or apathy?,9
post,3jurn7,2qh72,jokes,false,1441545920,https://old.reddit.com/r/Jokes/comments/3jurn7/pretty_good_one_liner/,self.jokes,,___________.,Pretty good one liner,4
post,3juq9t,2qh72,jokes,false,1441544978,https://old.reddit.com/r/Jokes/comments/3juq9t/a_redditor_has_sex_for_the_first_time/,self.jokes,https://www.reddit.com/r/Jokes/comments/3juq9t/a_redditor_has_sex_for_the_first_time/,,A Redditor has sex for the first time,1
post,3jupzu,2qh72,jokes,false,1441544775,https://old.reddit.com/r/Jokes/comments/3jupzu/intelligent_husband/,self.jokes,,[removed],Intelligent Husband,1
post,3juojk,2qh72,jokes,false,1441543765,https://old.reddit.com/r/Jokes/comments/3juojk/y_do_engineering_students_always_prefer_local/,self.jokes,,"The local author says;
“Jack &amp; Jill went up the hill to fetch a pail of water,
jack fell down and broke his crown and Jill came tumbling after""
&amp;
REFERENCE BOOK says;
“ 2 humans ascended a certain geological protuberance to collect
hydride of oxygen whose quantity is not specified.
One member Jack of rapid irregular disturbing movements encounter fatal logical gravitational error leading to complete disarray.
Other member whose scope lies within disarray descends down the geographical protuberance at an acceleration,
whose magnitude is controlled by the force of gravity.",Y do ENGINEERING students always prefer local author books then REFERENCE books..??,0
post,3juns4,2qh72,jokes,false,1441543172,https://old.reddit.com/r/Jokes/comments/3juns4/there_are_10_kinds_of_people/,self.jokes,,Those who get binary and those who don't.,There are 10 kinds of people.,0
post,3junny,2qh72,jokes,false,1441543093,https://old.reddit.com/r/Jokes/comments/3junny/polish_president_sends_a_telegram_to_the_german/,self.jokes,,[deleted],Polish president sends a telegram to the German Chancellor after the Soccer Game against Poland won by Germany last Friday,1
post,3jung3,2qh72,jokes,false,1441542924,https://old.reddit.com/r/Jokes/comments/3jung3/ambulances_are_the_original_transformers_because/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jung3/ambulances_are_the_original_transformers_because/,,Ambulances are the original Transformers because sometimes they transform mid-ride into hearses,0
post,3jundw,2qh72,jokes,false,1441542875,https://old.reddit.com/r/Jokes/comments/3jundw/do_you_know_the_difference_between_a_united/,self.jokes,,[deleted],Do you know the difference between a united states supreme court judge and an amature playwrite with dreams of hollywood?,1
post,3jun43,2qh72,jokes,false,1441542667,https://old.reddit.com/r/Jokes/comments/3jun43/i_was_going_to_tell_a_nirvana_joke_but/,self.jokes,,Nevermind.,"I was going to tell a Nirvana joke, but...",38
post,3jumvr,2qh72,jokes,false,1441542505,https://old.reddit.com/r/Jokes/comments/3jumvr/my_overweight_dad_has_been_running_9_miles_everday/,self.jokes,,[deleted],My overweight dad has been running 9 miles everday...,1
post,3jumpi,2qh72,jokes,false,1441542385,https://old.reddit.com/r/Jokes/comments/3jumpi/marines/,self.jokes,,"Two Marines boarded a quick shuttle flight out of Dallas, headed for Houston. One sat in the window seat, the other sat in the middle seat. Just before take-off, an Army soldier got on and took the aisle seat next to the two Marines. The Soldier kicked off his shoes, wiggled his toes and was settling in when the Marine in the window seat said, “I think I’ll get up and get a coke.” “No problem,” said the Soldier, “I’ll get it for you.” While he was gone, the Marine picked up the Soldier’s shoe and spit in it. When the Soldier returned with the coke, the Marine in the middle seat said, “That looks good, I think I’ll have one too.” Again, the Soldier obligingly went to fetch it and while he was gone, the Marine picked up the soldier’s other shoe and spit in it. The Soldier returned and they all sat back and enjoyed the rest of the short flight to Houston. As the plane was landing, the Soldier slipped his feet into his shoes and knew immediately what had happened. “How long must this go on?” the Soldier asked. “This fighting between our services? This hatred? This animosity? This spitting in shoes and peeing in cokes?”",Marines,2445
post,3jumem,2qh72,jokes,false,1441542161,https://old.reddit.com/r/Jokes/comments/3jumem/the_irish_mirror/,self.jokes,,[deleted],THE IRISH MIRROR,1325
post,3jum9a,2qh72,jokes,false,1441542049,https://old.reddit.com/r/Jokes/comments/3jum9a/puns_can_be_the_wurst_brat_i_sausage_you_might/,self.jokes,,[deleted],Puns can be the wurst. Brat I sausage you might appreciate this one.,0
post,3jum0e,2qh72,jokes,false,1441541875,https://old.reddit.com/r/Jokes/comments/3jum0e/i_refused_to_believe_my_roadworker_father_was/,self.jokes,,[deleted],I refused to believe my roadworker father was stealing from his job...,3
post,3julsu,2qh72,jokes,false,1441541694,https://old.reddit.com/r/Jokes/comments/3julsu/never_kiss_a_canary/,self.jokes,,"You'll get churpies! 
(It's a Canarial disease). ",Never kiss a Canary.,3
post,3julfn,2qh72,jokes,false,1441541400,https://old.reddit.com/r/Jokes/comments/3julfn/if_xmen_and_legend_of_korra_had_a_crossover_what/,self.jokes,,A Fassbender,If X-Men and Legend of Korra had a crossover what kind of bender would Magneto be?,1
post,3jul9q,2qh72,jokes,false,1441541285,https://old.reddit.com/r/Jokes/comments/3jul9q/how_does_a_syrian_family_have_a_meal/,self.jokes,,"The men provide the food and the women do the cooking, leaving the children to wash up afterwards. ",How does a Syrian family have a meal?,0
post,3jukb9,2qh72,jokes,false,1441540571,https://old.reddit.com/r/Jokes/comments/3jukb9/i_like_my_women_like_i_like_my_eggs/,self.jokes,,[deleted],I like my women like I like my eggs,0
post,3jujch,2qh72,jokes,false,1441539719,https://old.reddit.com/r/Jokes/comments/3jujch/what_do_you_call_the_continuous_urge_to_suck_dick/,self.jokes,,An addicktion,What do you call the continuous urge to suck dick?,2
post,3jujc3,2qh72,jokes,false,1441539710,https://old.reddit.com/r/Jokes/comments/3jujc3/long_winded_so_the_local_church_bell_ringer_dies/,self.jokes,,"There is a small village in rural England, which has a church. In the church lives a priest and the bell ringer. One morning the priest doesn't hear the morning bell ring so he goes to the bell ringers room to check on him. When he enters the room he sees the bell ringer dead in his bed.

The priest, although he is upset, makes some flyers about new bell ringer auditions and sticks them to every lamp-post in the village. The next day there is a huge line of people queuing outside the Church. The priest, surprised by the amount of people, eagerly welcomes them in one by one to see who is the best ringer. Around 200 people try out and the line slowly gets shorter and shorter until everyone has tried to impress the priest with their bell ringing. 

Although there were some brilliant ringers that day non of them were up to the standards of the old bell ringer. The priest slumped in his chair, disappointed with the days outcome when suddenly he hears a bang on the door. He opens the door and doesn't see anyone..

""Down here!"" A man shouts. The priest looks down and before him stood a man with no arms or legs. ""I hope I'm not late for the bell ringing try outs"" the man said.

""err... no you're not, come this way"" the priest said unsurely. He carried the man up to the bell tower and placed him in front of the bell and the rope to ring it. The man starred at he bell for a while until he began to hit his head on it.. hard.. again.. and again. The priest was in complete awe at his amazing skills. 

The man carried on.. hitting his head on the bell harder and harder, fastest and faster. Blood begins to appear.. trickling down his face but he keeps on going... eventually he falls to the ground. The priest kneels down to inspect him... he is unconscious.

The priest immediately runs into the village to go and get help. ""Help! Somebody help!"" he shouted. He gathered a small crowd of people and took them to church. They all gathered around the unconscious man. Upon closer inspection they realise he was dead.. the priest begins to cry.. ""He was brilliant.. the best I have ever heard.... I didn't even know his name! Who was this man!?""

The crowd look at each other until one man stood out and said:

""I don't know his name.. but his face rings a bell.""",[Long Winded] So the local church bell ringer dies.,25
post,3juj8k,2qh72,jokes,false,1441539633,https://old.reddit.com/r/Jokes/comments/3juj8k/how_many_germans_does_it_take_to_screw_in_a/,self.jokes,,One. They are efficient and not very funny.,How many germans does it take to screw in a lightbulb?,0
post,3jui5w,2qh72,jokes,false,1441538705,https://old.reddit.com/r/Jokes/comments/3jui5w/what_is_the_difference_between_a_chair_and_a_cock/,self.jokes,,Be careful where you sit down,What is the difference between a chair and a cock?,0
post,3jui4y,2qh72,jokes,false,1441538687,https://old.reddit.com/r/Jokes/comments/3jui4y/i_put_my_grandma_on_speed_dial/,self.jokes,,"Instagram is a thing, right? ",I put my grandma on speed dial.,0
post,3juhel,2qh72,jokes,false,1441538035,https://old.reddit.com/r/Jokes/comments/3juhel/someone_stole_my_coffee/,self.jokes,,He was charged with mugging. ,Someone stole my coffee.,136
post,3juhd9,2qh72,jokes,false,1441538003,https://old.reddit.com/r/Jokes/comments/3juhd9/i_was_just_watching_the_chinese_parade_i_was/,self.jokes,,[deleted],I was just watching the Chinese parade I was impressed.....,0
post,3jugqn,2qh72,jokes,false,1441537433,https://old.reddit.com/r/Jokes/comments/3jugqn/the_other_day_a_clown_held_the_door_open_for_me/,self.jokes,,It was a nice jester. ,"The other day, a clown held the door open for me.",8
post,3jugf2,2qh72,jokes,false,1441537115,https://old.reddit.com/r/Jokes/comments/3jugf2/buddha_is_not_a_god/,self.jokes,,But he sure looks like he ate one,Buddha is not a god,0
post,3jug4r,2qh72,jokes,false,1441536829,https://old.reddit.com/r/Jokes/comments/3jug4r/whats_white_and_wears_red_checked_trousers/,self.jokes,,Rupert the fridge.,What's white and wears red checked trousers....,2
post,3jufre,2qh72,jokes,false,1441536472,https://old.reddit.com/r/Jokes/comments/3jufre/100m_dash/,self.jokes,,"A girl says to her friend ""The last time I had sex was like the 100 meter dash""

Her friend says ""What, over in 6 seconds?""

""No, with 8 black men and a gun.""",100m Dash,5841
post,3jufd1,2qh72,jokes,false,1441536125,https://old.reddit.com/r/Jokes/comments/3jufd1/i_saw_a_weird_competition_yesterday_the_first/,self.jokes,,So I entered myself.,I saw a weird competition yesterday - The first person to successfully have intercourse with them self wins.,52
post,3juf4f,2qh72,jokes,false,1441535887,https://old.reddit.com/r/Jokes/comments/3juf4f/op/,self.jokes,https://www.reddit.com/r/Jokes/comments/3juf4f/op/,,OP,0
post,3juemt,2qh72,jokes,false,1441535421,https://old.reddit.com/r/Jokes/comments/3juemt/what_do_you_say_when_a_robot_explodes_into_pieces/,self.jokes,,Rest in pieces. I'll show myself out now.,What do you say when a robot explodes into pieces?,2
post,3juedt,2qh72,jokes,false,1441535157,https://old.reddit.com/r/Jokes/comments/3juedt/so_a_man_walks_into_a_bar/,self.jokes,,[deleted],So a man walks into a bar,0
post,3jue4s,2qh72,jokes,false,1441534941,https://old.reddit.com/r/Jokes/comments/3jue4s/01021183715_부산출장안마부산출장마사지부산출장아가씨부산_전지역/,self.jokes,,[removed],"010-2118-3715 부산출장안마,부산출장마사지,부산출장아가씨,부산 전지역 출장안마,마사지,서비스,업소,업체,모텔바리,아가씨,걸,녀,유흥,방문,콜걸",1
post,3judww,2qh72,jokes,false,1441534748,https://old.reddit.com/r/Jokes/comments/3judww/oc_what_did_the_auditors_say_to_the_south/,self.jokes,,"Hello, I'm here to Peru-se your inventory.",(OC) What did the auditors say to the South American shopkeeper?,1
post,3judr4,2qh72,jokes,false,1441534616,https://old.reddit.com/r/Jokes/comments/3judr4/so_a_man_dies_and_is_neither_good_or_bad/,self.jokes,,[deleted],"So a man dies, and is neither good or bad.",0
post,3judqq,2qh72,jokes,false,1441534609,https://old.reddit.com/r/Jokes/comments/3judqq/an_englishman_an_irishman_and_a_scotsman/,self.jokes,,"An Englishman, an Irishman, and a Scotsman were all builders sitting at the top of their current construction site for lunch. The Englishman opened his sandwich and turned to the others to say: 
""Bloody hell I've got Ham and Cheese again!""
The Irishman looks at his sandwich and says: ""Aye, I have tuna sandwiches yet again!"". 
Likewise, the Scotsman commented on his lunch: ""I've got egg as always!""

The three men exchanged looks before the Englishman decided: ""I've had enough of this! If I end up with Ham and Cheese again I'm going to jump off this building!!"" The other two nodded in agreement stating that they would too.

The next day the Englishman had ham and cheese, the Irishman had tuna, and the Scotsman had egg. And, as promised the day before, they jumped off the building.


At their funeral a week later, their wives, sobbing, began to talk. 
The Englishman's wife said ""If only he had told me that he didn't like Ham and Cheese I would've made him something else!!"" 
The Irishman's wife agreed ""I didn't know that he hated tuna!"" 
Then the Scotsman's wife turned around and said ""I don't know what you're on about - he made his own bloody lunch!""","An Englishman, an Irishman, and a Scotsman...",4
post,3judo7,2qh72,jokes,false,1441534547,https://old.reddit.com/r/Jokes/comments/3judo7/pet_diaries/,self.jokes,,"Excerpts from a Dog's Diary:

* 8:00 am - Dog food! My favourite thing!
* 9:30 am - A car ride! My favourite thing!
* 9:40 am - A walk in the park! My favourite thing!
* 10:30 am - Got rubbed and petted! My favourite thing!
* 12:00 pm - Lunch! My favourite thing!
* 1:00 pm - Played in the yard! My favourite thing!
* 3:00 pm - Wagged my tail! My favourite thing!
* 5:00 pm - Milk bones! My favourite thing!
* 7:00 pm - Got to play ball! My favourite thing!
* 8:00 pm - Wow! Watched TV with the people! My favourite thing!
* 11:00 pm - Sleeping on the bed! My favourite thing!

Excerpts from a Cat's Diary:

Day 983 of my captivity.

My captors continue to taunt me with bizarre little dangling objects. They dine lavishly on fresh meat, while the other inmates and I are fed hash or some sort of dry nuggets. Although I make my contempt for the rations perfectly clear, I nevertheless must eat something in order to keep up my strength. The only thing that keeps me going is my dream of escape. In an attempt to disgust them, I once again vomit on the carpet. 
Today I decapitated a mouse and dropped its headless body at their feet. I had hoped this would strike fear into their hearts, since it clearly demonstrates what I am capable of. However, they merely made condescending comments about what a ""good little hunter"" I am.

Bastards!

There was some sort of assembly of their accomplices tonight. I was placed in solitary confinement for the duration of the event. However, I could hear the noises and smell the food. I overheard that my confinement was due to the power of ""allergies."" I must learn what this means, and how to use it to my advantage.

Today I was almost successful in an attempt to assassinate one of my tormentors by weaving around his feet as he was walking. I must try this again tomorrow - but at the top of the stairs. 

I am convinced that the other prisoners here are flunkies and snitches. The dog receives special privileges. He is regularly released - and seems to be more than willing to return. He is obviously retarded. The bird has got to be an informant. I observe him communicate with the guards regularly. I am certain that he reports my every move. My captors have arranged protective custody for him in an elevated cell, so he is safe. For now...",Pet Diaries:,106
post,3judnx,2qh72,jokes,false,1441534542,https://old.reddit.com/r/Jokes/comments/3judnx/the_old_joke_i_assume_this_site_was_named_after_a/,self.jokes,,[deleted],The old joke I assume this site was named after - A chicken walks into a library...,78
post,3jucwb,2qh72,jokes,false,1441533832,https://old.reddit.com/r/Jokes/comments/3jucwb/rich_man/,self.jokes,,"A wealthy man was driving in his car when he saw two men along the roadside eating grass.
Disturbed by the sight, he ordered his driver to stop and he got out to investigate. He asked one man, ""Why are you eating grass?""
""We don't have any money for food,"" the poor man replied.
""We have to eat grass.""
""Well, then, you can come with me to my house and I'll feed you,"" the man said.
""But sir, I have a wife and five children with me. They are over there, under that tree"".
""Bring them along,"" the rich man replied. Turning to the other poor man he stated, ""You come with us, too.""
The second man, in a pitiful voice then said, ""But sir, I also have a wife and seven children with me!""
""Bring them all, as well,"" the man answered. They all entered the car, which was no easy task, even for a car as large as it was.
One of the poor fellows turned to the rich man and said, ""Sir, you are too kind. Thank you for taking all of us with you.""
The manager replied, ""Glad to do it. You'll really love my place; the grass is almost 1 meter high!""",Rich Man,0
post,3jucm5,2qh72,jokes,false,1441533548,https://old.reddit.com/r/Jokes/comments/3jucm5/why_do_bees_hum/,self.jokes,,Because they can't remember the lyrics,Why do bees hum?,4
post,3jucem,2qh72,jokes,false,1441533327,https://old.reddit.com/r/Jokes/comments/3jucem/a_man_who_says_his_wife_cannot_take_a_joke/,self.jokes,,[deleted],A man who says his wife cannot take a joke...,1
post,3jubhj,2qh72,jokes,false,1441532412,https://old.reddit.com/r/Jokes/comments/3jubhj/fishes/,self.jokes,,What does a fish say when it hits a concrete wall? ,Fishes.,1
post,3jubh5,2qh72,jokes,false,1441532404,https://old.reddit.com/r/Jokes/comments/3jubh5/i_have_two_friends_who_always_compete_against/,self.jokes,,But they always end in a draw,I have two friends who always compete against each other in art competitions,26
post,3jubem,2qh72,jokes,false,1441532335,https://old.reddit.com/r/Jokes/comments/3jubem/mum_where_do_i_hang_the_clothes_the_hanging_lines/,self.jokes,,"Son, just hang them in the gallows. No one would know.","Mum, where do I hang the clothes. The hanging line's gone.",2
post,3jub6v,2qh72,jokes,false,1441532141,https://old.reddit.com/r/Jokes/comments/3jub6v/bridge_is_like_sex/,self.jokes,,"If you don't have a good partner, you'd better have a good hand.",Bridge is like sex,4
post,3juaud,2qh72,jokes,false,1441531802,https://old.reddit.com/r/Jokes/comments/3juaud/my_muslim_friends/,self.jokes,,"So I've got a pretty diverse friend group, of which includes several Muslims.

There's:

•That guy who lives between two other houses- Ali

•That guy with a sausage in his hair - Hamed

•Oh and that other guy, who looks like he has two sausages in his hair! Mohammed!

Bonus :(《hint》May require some punjabi). That guy with a receding hairline -Ikbal


No religious hate intended ♡♥",My Muslim friends,0
post,3juamq,2qh72,jokes,false,1441531593,https://old.reddit.com/r/Jokes/comments/3juamq/pass_me_the_hammafor/,self.jokes,https://www.reddit.com/r/Jokes/comments/3juamq/pass_me_the_hammafor/,,Pass me the hamma-for,0
post,3jua0l,2qh72,jokes,false,1441530988,https://old.reddit.com/r/Jokes/comments/3jua0l/johnny_and_the_cow_short_and_sweet/,self.jokes,,"I heard a tale once about a boy  called Johnny. He impressed his whole village by his unique ability to sit for hours underneath a cow.

He was rewarded with a pat on the head.",Johnny and the cow - short and sweet,2
post,3jua0h,2qh72,jokes,false,1441530987,https://old.reddit.com/r/Jokes/comments/3jua0h/updatekentucky_vs_south_carolina_live_online/,self.jokes,,[removed],Update:Kentucky vs South Carolina live online,1
post,3ju9rr,2qh72,jokes,false,1441530783,https://old.reddit.com/r/Jokes/comments/3ju9rr/if_a_man_says_hes_going_to_fix_it_he_is_going_to/,self.jokes,,[deleted],"If a man says he's going to fix it, he IS going to fix it.",0
post,3ju8hn,2qh72,jokes,false,1441529497,https://old.reddit.com/r/Jokes/comments/3ju8hn/good_answer/,self.jokes,,"A white couple gets a black child.
Angry husband asks- You white, Me white. Why is baby black?
Wife- You hot, Me hot. Baby burnt!

",Good Answer,1
post,3ju6o1,2qh72,jokes,false,1441527744,https://old.reddit.com/r/Jokes/comments/3ju6o1/special_occasions/,self.jokes,,"Once when I was little and had just started to learn to read, I went to the bathroom and noticed a box with the word ""napkins"" on it.
I was proud that I could read that word but puzzled and asked my mom a why she was keeping ""napkins"" in the bathroom. 
Didn't they belong in the kitchen?

Not wanting to burden me with unnecessary facts, she told me that they were for ""special occasions"".

A few months later - it's Thanksgiving, and Mom had assignments for all of us.

Mine was to set the table.

Now the fun started.
When the guests arrived, my uncle came in first and immediately burst into laughter. 
Next came his wife who gasped,and then giggled.
Then came my father, who roared with laughter.

Then came mom, who almost died of embarrassment when she saw each place setting on the table with a Kotex napkin at each plate, with the fork carefully arranged on top. I had even tucked in the wings!

My mother asked me why I used these and, of course, my response sent the other adults into further fits of laughter.

""But, Mom, you said that they were for special occasions!""",Special Occasions,0
post,3ju49r,2qh72,jokes,false,1441525661,https://old.reddit.com/r/Jokes/comments/3ju49r/whats_the_worst_last_words_your_exgf_can_say_to/,self.jokes,,"""I do."" ",What's the worst last words your EX-GF can say to you?,16
post,3ju3nt,2qh72,jokes,false,1441525106,https://old.reddit.com/r/Jokes/comments/3ju3nt/a_chicken_and_an_egg_lie_together_in_bed/,self.jokes,,[deleted],A chicken and an egg lie together in bed,0
post,3ju3cp,2qh72,jokes,false,1441524827,https://old.reddit.com/r/Jokes/comments/3ju3cp/yesterday_i_took_my_grandchildren_to_the_park_a/,self.jokes,,"I was outraged,

her kids weren't even hot.","Yesterday I took my grandchildren to the park, a Woman came up to me and accused me of being a paedophile.",3
post,3ju2qx,2qh72,jokes,false,1441524330,https://old.reddit.com/r/Jokes/comments/3ju2qx/what_is_empty_and_spins_round_and_round/,self.jokes,,A Malaysian Airlines baggage claim. ,What is empty and spins round and round?,34
post,3ju2ac,2qh72,jokes,false,1441523995,https://old.reddit.com/r/Jokes/comments/3ju2ac/mr_president_two_brazilian_soldiers_were_executed/,self.jokes,,[deleted],"""Mr. President, two Brazilian soldiers were executed yesterday in Iraq.""",0
post,3ju20f,2qh72,jokes,false,1441523751,https://old.reddit.com/r/Jokes/comments/3ju20f/what_did_adolf_hitler_get_his_niece_for_her/,self.jokes,,"An easy bake oven.

i don't give two shits if you heard this before or if this is a repost, this is mainly for shits and giggles =)",What did Adolf Hitler get his niece for her birthday?,0
post,3ju1xl,2qh72,jokes,false,1441523686,https://old.reddit.com/r/Jokes/comments/3ju1xl/i_identify_as_a_sexual_atheist/,self.jokes,,I dont believe I'll ever get laid. ,I identify as a Sexual Atheist,4
post,3ju1k0,2qh72,jokes,false,1441523317,https://old.reddit.com/r/Jokes/comments/3ju1k0/a_jewish_kid_asks_his_father_for_twenty_dollars/,self.jokes,,"His father replied, ""ten dollars, what in the world do you need five dollars for, I'd be happy to give you a dollar, here's one cent."" ",A Jewish kid asks his father for twenty dollars.,0
post,3ju1bp,2qh72,jokes,false,1441523095,https://old.reddit.com/r/Jokes/comments/3ju1bp/806_mr_president_two_brazilian_soldiers_were/,self.jokes,,[deleted],"806 ""Mr. President, two Brazilian soldiers were executed yesterday in Iraq.""",1
post,3ju185,2qh72,jokes,false,1441522985,https://old.reddit.com/r/Jokes/comments/3ju185/the_european_commission_has_just_announced_an/,self.jokes,,"...whereby English will be the official language of the European Union rather than German, which was the other possibility.
As part of the negotiations, the British Government conceded that English spelling had some room for improvement and has accepted a 5- year phase-in plan that would become known as ""Euro-English"".
In the first year, ""s"" will replace the soft ""c"". Sertainly, this will make the sivil servants jump with joy. The hard ""c"" will be dropped in favour of ""k"". This should klear up konfusion, and keyboards kan have one less letter.
There will be growing publik enthusiasm in the sekond year when the troublesome ""ph"" will be replaced with ""f"". This will make words like fotograf 20% shorter.
In the 3rd year, publik akseptanse of the new spelling kan be expekted to reach the stage where more komplikated changes are possible. Governments will enkourage the removal of double letters which have always ben a deterent to akurate speling. Also, al wil agre that the horibl mes of the silent ""e"" in the languag is disgrasful and it should go away.
By the 4th yer people wil be reseptiv to steps such as replasing ""th"" with ""z"" and ""w"" with ""v"".
During ze fifz yer, ze unesesary ""o"" kan be dropd from vords kontaining ""ou"" and after ziz fifz yer, ve vil hav a reil sensi bl riten styl.
Zer vil be no mor trubl or difikultis and evrivun vil find it ezi tu understand ech oza. Ze drem of a united urop vil finali kum tru!
Und efter ze fifz yer, ve vil al be speking German like zey vunted in ze forst plas.",The European Commission has just announced an agreement,0
post,3ju123,2qh72,jokes,false,1441522829,https://old.reddit.com/r/Jokes/comments/3ju123/what_do_you_call_75_year_old_john_cena/,self.jokes,,John Cenile.,What do you call 75 year old John Cena?,12
post,3ju0vt,2qh72,jokes,false,1441522657,https://old.reddit.com/r/Jokes/comments/3ju0vt/watch_college_football_live_online/,self.jokes,,[removed],WATCH COLLEGE FOOTBALL LIVE ONLINE,0
post,3ju0ux,2qh72,jokes,false,1441522626,https://old.reddit.com/r/Jokes/comments/3ju0ux/how_do_you_fit_15_jews_into_a_car/,self.jokes,,"2 in the front,3 in the back,and the rest in the ash tray.",How do you fit 15 Jews into a car?,1
post,3ju0tu,2qh72,jokes,false,1441522601,https://old.reddit.com/r/Jokes/comments/3ju0tu/what_do_you_get_when_you_cross_a_joke_with_a/,self.jokes,https://www.reddit.com/r/Jokes/comments/3ju0tu/what_do_you_get_when_you_cross_a_joke_with_a/,,What do you get when you cross a joke with a rhetorical question?,22
post,3ju0r9,2qh72,jokes,false,1441522546,https://old.reddit.com/r/Jokes/comments/3ju0r9/how_much_does_the_turtle_cross_the_free_way_old/,self.jokes,,"Mary, Mother of Jesus, is trying to pull a bullfrog out of his wife's vagina. An old man lives in a retirement home and realizes that he has lost 10 lbs. as promised. On July 4, 3055, Steel revealed a massive construct the size of a submarine.You can do all the work and the fat guy with the orange head, introduces himself, and offers to buy the bullfrog for $100,000.",How much does the turtle cross the free way? old man's advice,0
post,3ju0av,2qh72,jokes,false,1441522076,https://old.reddit.com/r/Jokes/comments/3ju0av/poland_is_so_obscene/,self.jokes,,[deleted],Poland is so obscene...,1
post,3ju0a0,2qh72,jokes,false,1441522049,https://old.reddit.com/r/Jokes/comments/3ju0a0/whats_the_difference_between_a_jew_and_a_pizza/,self.jokes,,A pizza doesn't scream when you put it in the oven.,What's the difference between a jew and a pizza?,0
post,3ju054,2qh72,jokes,false,1441521937,https://old.reddit.com/r/Jokes/comments/3ju054/the_dead_batteries_were_given_out_to_people/,self.jokes,,[deleted],The dead batteries were given out to people...,2
post,3ju04n,2qh72,jokes,false,1441521925,https://old.reddit.com/r/Jokes/comments/3ju04n/a_new_zealander_visits_us/,self.jokes,,"A New Zealander lands in NYC. His American friend comes to pick him at JFK. American friend asks, where do you want to visit first? NZer says, rocky mountain national park in Colorado. His American friend is real surprised. Why not visit Manhattan or California or Florida first? Why do you want to visit Colorado first? I mean it is real nice place, but why?

NZer says, I want to have wild sex.

PS: original joke. If no one understands, I can perhaps provide a clue",A New Zealander visits US,0
post,3ju003,2qh72,jokes,false,1441521817,https://old.reddit.com/r/Jokes/comments/3ju003/most_guys_experiment_with_homosexuality_in_college/,self.jokes,,I experimented in Sunday School,Most guys experiment with homosexuality in college...,1
post,3jtzgi,2qh72,jokes,false,1441521351,https://old.reddit.com/r/Jokes/comments/3jtzgi/there_are_two_types_of_people_in_the_world/,self.jokes,,"...those who pee in the shower, and liars.",There are two types of people in the world...,17
post,3jtzfg,2qh72,jokes,false,1441521323,https://old.reddit.com/r/Jokes/comments/3jtzfg/a_black_jewish_boy_runs_home_from_school_one_day/,self.jokes,," ...and asks his father, “Daddy, am I more Jewish or more black?”  The dad replies, “Why do you want to know, son?” “Because a kid at school is selling a bike for $50 and I want to know if I should talk him down to $40 or just steal it!”",A black Jewish boy runs home from school one day...,159
post,3jtza0,2qh72,jokes,false,1441521204,https://old.reddit.com/r/Jokes/comments/3jtza0/whats_the_closest_synonym_to_a_love_boat/,self.jokes,,A relation-ship.,What's the closest synonym to a love boat?,6
post,3jtyt8,2qh72,jokes,false,1441520852,https://old.reddit.com/r/Jokes/comments/3jtyt8/a_christian_a_buddhist_an_atheist_and_an_agnostic/,self.jokes,,"All of a sudden, the plane is about to crash, and so the passengers need to jump off due to the lack of parachutes.

The Christian jumps off first and says, ""God will save me!"" and God saves him.

The Buddhist then jumps off and says, ""Buddha will save me!"" and Buddha saves him.

Now because the atheist didn't believe in any higher being, he says, ""Nobody will save me!"" So nobody saves him and he dies.

The agnostic then says to himself, ""Wow, what an idiot."" So he decides to become Buddhist temporarily, as he did not reject the idea of a God as an agnostic. He jumps off and says, ""Buddha will save me!"" and Buddha saves him in midair. 

Then he said, ""Thank God that worked."" Buddha then drops him and he dies.","A Christian, a Buddhist, an atheist, and an agnostic are on a plane",15
post,3jtwyg,2qh72,jokes,false,1441519392,https://old.reddit.com/r/Jokes/comments/3jtwyg/pakistani_chat_rooms_online_without_registration/,self.jokes,,[removed],Pakistani Chat Rooms Online Without Registration,0
post,3jtw0h,2qh72,jokes,false,1441518586,https://old.reddit.com/r/Jokes/comments/3jtw0h/what_did_the_old_billy_bobs_eat_at_mcdonalds/,self.jokes,,McChicken-killer... Yeah I'm really stoned smoked a chicken killer and ate McDonald's,What did the old billy bobs eat at McDonald's?,0
post,3jtvh1,2qh72,jokes,false,1441518130,https://old.reddit.com/r/Jokes/comments/3jtvh1/ill_bet_that_referees_are_especially_in_favor_of/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jtvh1/ill_bet_that_referees_are_especially_in_favor_of/,,I'll bet that referees are especially in favor of whistleblower protection laws.,0
post,3jturq,2qh72,jokes,false,1441517600,https://old.reddit.com/r/Jokes/comments/3jturq/two_elderly_couples_were_enjoying_friendly/,self.jokes,,"Two elderly couples were enjoying friendly conversation when... one of the men asked the other, ""Fred, how was the memory clinic you went to last month?""

""Outstanding,"" Fred replied. ""They taught us all the latest psychological techiniques-visulization, association-it made a huge difference for me.""

""That's great! What was the name of the clinic?""

Fred went blank He thought and thought, but couldn't remember.

Then a smile broke across his face and he asked, ""What do you call that flower with the long stem and thorns?""

""You mean a rose?""

""Yes, that's it!"" He turned to his wife. . .""Rose, what was the name of that clinic?""

(copied from http://www.ahajokes.com/age49.html)",Two elderly couples were enjoying friendly conversation when...,4
post,3jtulu,2qh72,jokes,false,1441517498,https://old.reddit.com/r/Jokes/comments/3jtulu/why_do_white_girls_only_travel_in_packs_of_3s/,self.jokes,,Because omg they can't even.,Why do white girls only travel in packs of 3's?,1
post,3jttjo,2qh72,jokes,false,1441516747,https://old.reddit.com/r/Jokes/comments/3jttjo/whats_the_difference_between_a_chickpea_and_a/,self.jokes,,I've never had a garbanzo bean on my chest. ,What's the difference between a chickpea and a garbanzo bean...?,13
post,3jtt6x,2qh72,jokes,false,1441516509,https://old.reddit.com/r/Jokes/comments/3jtt6x/kanye_west_announced_that_he_was_going_to_run_for/,self.jokes,,[deleted],Kanye West announced that he was going to run for president in 2020,0
post,3jtt57,2qh72,jokes,false,1441516473,https://old.reddit.com/r/Jokes/comments/3jtt57/a_man_walks_into_a_bar/,self.jokes,,His friends ducked.,A man walks into a bar...,0
post,3jtsz9,2qh72,jokes,false,1441516365,https://old.reddit.com/r/Jokes/comments/3jtsz9/i_exercise_religiously/,self.jokes,,I go to the gym for an hour on Sunday morning and then don't think about it again for the rest of the week.,I exercise religiously,237
post,3jtsmr,2qh72,jokes,false,1441516103,https://old.reddit.com/r/Jokes/comments/3jtsmr/whats_the_difference_between_a_mechanical_and_a/,self.jokes,,One builds weapons and the other build targets. ,What's the difference between a mechanical and a civil engineer?,150
post,3jtsad,2qh72,jokes,false,1441515880,https://old.reddit.com/r/Jokes/comments/3jtsad/a_guy_named_michael_was_rushed_to_the_emergency/,self.jokes,,I guess you could say it was open Mike night.,A guy named Michael was rushed to the emergency room one night and had to have heart surgery..,2
post,3jtrnw,2qh72,jokes,false,1441515449,https://old.reddit.com/r/Jokes/comments/3jtrnw/why_do_sorority_girls_travel_in_packs_of_1_3_5_or/,self.jokes,,Because they can't even.,"Why Do Sorority Girls Travel In Packs Of 1, 3, 5 or 7?",6
post,3jtr6r,2qh72,jokes,false,1441515088,https://old.reddit.com/r/Jokes/comments/3jtr6r/i_was_talking_with_my_lunkheads_boyfriend_the/,self.jokes,,"And I told him about my new research. I'm a biologist studying primate reproductive organs, and we are doing new research on a substance produced in urine by certain lemurs called nisch. It's essentially an acid designed to keep predators away, but it hurts like hell to pass it. 

I mentioned to him that I'm glad I'm not a lemur, 
because  that shit burns. ""I'm eternally thankful thank I can't pee nisch""

""Wait, what? I had no idea you were a lesbian!""",I was talking with my lunkheads boyfriend the other day,0
post,3jtqjt,2qh72,jokes,false,1441514674,https://old.reddit.com/r/Jokes/comments/3jtqjt/little_johnny_is_in_his_bedroom_when_his_mother/,self.jokes,,"She says to him, ""Little Johnny, we're going to the neighbor's house tonight for dinner to celebrate the birth of their new baby.""

""Okay, mommy,"" he replies.

""Now listen carefully: the baby was born without ears. I don't want you making ear jokes or hearing jokes or anything of the sort. If you do, you'll be grounded for a month!""

""Okay, mommy,"" Little Johnny says.

They go to the neighbor's house and have a lovely 3-course meal. After dessert is cleared away, they all go into the nursery to see the baby, sleeping soundly in his bassinet.

Little Johnny is peeking up over the side in obvious fascination. The baby's mother smiles down at Johnny and says, ""What do you think of the baby, Johnny?""

""Oh, ma'am, that is a beautiful baby! He has such beautiful hands and beautiful feet and beautiful eyes. Does he see okay?""

""He sure does,"" she says with a bright smile, ""The doctor says he's be blessed with perfect 20/20 vision.""

""That's good because if he needed glasses, he'd be fucked.""",Little Johnny Is In His Bedroom When His Mother Walks In,7
post,3jtpy4,2qh72,jokes,false,1441514285,https://old.reddit.com/r/Jokes/comments/3jtpy4/a_man_boarded_an_airplane_and_took_his_seat_as_he/,self.jokes,,[deleted],"A man boarded an airplane and took his seat. As he settled in, he glanced Up and saw the most beautiful woman boarding the plane",0
post,3jtps4,2qh72,jokes,false,1441514162,https://old.reddit.com/r/Jokes/comments/3jtps4/why_did_the_teacher_cross_her_eyes/,self.jokes,,Because she couldn't control her pupils.,Why did the teacher cross her eyes?,6
post,3jtpru,2qh72,jokes,false,1441514158,https://old.reddit.com/r/Jokes/comments/3jtpru/did_you_guys_know_that_water_can_talk/,self.jokes,,Water you talking about?,Did you guys know that water can talk?,2
post,3jtopn,2qh72,jokes,false,1441513454,https://old.reddit.com/r/Jokes/comments/3jtopn/whats_a_bears_favorite_paint_company/,self.jokes,,[deleted],What's a bear's favorite paint company?,0
post,3jtodt,2qh72,jokes,false,1441513250,https://old.reddit.com/r/Jokes/comments/3jtodt/what_do_you_call_fake_spaghetti/,self.jokes,,An impasta!,What Do You Call Fake Spaghetti?,1
post,3jtobm,2qh72,jokes,false,1441513205,https://old.reddit.com/r/Jokes/comments/3jtobm/a_man_boarded_an_airplane_and_took_his_seat/,self.jokes,,[deleted],A man boarded an airplane and took his seat.,6
post,3jto4t,2qh72,jokes,false,1441513081,https://old.reddit.com/r/Jokes/comments/3jto4t/did_you_hear_about_the_guy_who_ate_his_trousers/,self.jokes,,He pooped his pants!,Did you hear about the guy who ate his trousers?,29
post,3jtnoa,2qh72,jokes,false,1441512779,https://old.reddit.com/r/Jokes/comments/3jtnoa/americas_a_terrorist_country_why/,self.jokes,,[removed],"America's a terrorist country, why?",0
post,3jtno8,2qh72,jokes,false,1441512778,https://old.reddit.com/r/Jokes/comments/3jtno8/whats_the_difference_between_a_piano_and_tuna/,self.jokes,,You can tuna piano but you can't tuna fish.,What's the difference between a piano and tuna?,0
post,3jtnbc,2qh72,jokes,false,1441512569,https://old.reddit.com/r/Jokes/comments/3jtnbc/these_two_kids_want_to_be_roasted/,self.jokes,,[removed],These two kids want to be roasted!,0
post,3jtn42,2qh72,jokes,false,1441512450,https://old.reddit.com/r/Jokes/comments/3jtn42/jared_from_subway_ended_his_career_the_same_way/,self.jokes,,Trying to get into small pants.,Jared from Subway ended his career the same way he started it.,3
post,3jtmmg,2qh72,jokes,false,1441512178,https://old.reddit.com/r/Jokes/comments/3jtmmg/two_sperms_are_talking_with_each_other/,self.jokes,,"""Hey man, how long till we get the ovaries?""

""Long way still, we just passed the throat.""",Two sperms are talking with each other...,20
post,3jtmlb,2qh72,jokes,false,1441512159,https://old.reddit.com/r/Jokes/comments/3jtmlb/when_homer_simpson_plays_dungeons_dragons/,self.jokes,,He uses a D'oh!-decahedron.,When Homer Simpson plays Dungeons &amp; Dragons...,1
post,3jtmkb,2qh72,jokes,false,1441512141,https://old.reddit.com/r/Jokes/comments/3jtmkb/a_man_boarded_an_airplane_and_took_his_seat_as_he/,self.jokes,,"The most beautiful woman boarding the plane. He soon realized She was heading straight towards his seat. As fate would have it, she took The seat right beside his. Eager to strike up a conversation he blurted out, “Business trip or pleasure?”
She turned, smiled and said, “Business. I’m going to the Annual Nymphomaniacs of America Convention in Boston.""
He swallowed hard. Here was the most gorgeous woman he had ever seen Sitting next to him, and she was going to a meeting of nymphomaniacs!
Struggling to maintain his composure, he calmly asked, “What’s your Business at this convention?”
“Lecturer,” she responded. “I use information that I have learned from my Personal experiences to debunk some of the popular myths about sexuality.”
“Really?” he said. “And what kind of myths are there?”
“Well,” she explained, “one popular myth is that African-American men are The most well-endowed of all men, when in fact it is the Native American Indian who is most likely to possess that trait. Another popular myth is That Frenchmen are the best lovers, when actually it is men of Mexican Descent who are the best. I have also discovered that the lover with Absolutely the best stamina is the Southern Redneck.”
Suddenly the woman became a little uncomfortable and blushed.. “I’m Sorry,” she said, “I shouldn't really be discussing all of this with you. I don’t Even know your name.”
“Tonto,” the man said, “Tonto Gonzales, but my friends call me Bubba"".","A man boarded an airplane and took his seat. As he settled in, he glanced Up and saw",0
post,3jtmfg,2qh72,jokes,false,1441512064,https://old.reddit.com/r/Jokes/comments/3jtmfg/knock_knockwhos_theremaijumaiju_who/,self.jokes,,[deleted],"""Knock Knock"",""Who's there?"",""Maiju"",""Maiju who?""",0
post,3jtlz4,2qh72,jokes,false,1441511778,https://old.reddit.com/r/Jokes/comments/3jtlz4/when_i_die_i_want_to_be_buried_by_my_group_members/,self.jokes,,..so they can let me down one last time.,When I die I want to be buried by my group members...,0
post,3jtln9,2qh72,jokes,false,1441511575,https://old.reddit.com/r/Jokes/comments/3jtln9/what_do_you_call_it_when_bob_dylan_sucks_your/,self.jokes,,The answer my friend... is blowing in the wind. The answer is blowing in the wind.,What do you call it when Bob Dylan sucks your dick in a hurricane?,12
post,3jtl9r,2qh72,jokes,false,1441511332,https://old.reddit.com/r/Jokes/comments/3jtl9r/an_illinois_man_left_the_cold_streets_of_chicago/,self.jokes,,[deleted],An Illinois man left the cold streets of Chicago for a vacation in Florida.,16
post,3jtl8i,2qh72,jokes,false,1441511309,https://old.reddit.com/r/Jokes/comments/3jtl8i/my_friend_just_said_this/,self.jokes,,Never be a half assed dog owner... It'll bite you in the ass every time,My friend just said this:,0
post,3jtkri,2qh72,jokes,false,1441511011,https://old.reddit.com/r/Jokes/comments/3jtkri/what_is_in_common_between_a_napkin_and_a_person/,self.jokes,,"If you sleep with a person, he/she is ur nap-kin.",What is in common between a napkin and a person?,0
post,3jtjwk,2qh72,jokes,false,1441510486,https://old.reddit.com/r/Jokes/comments/3jtjwk/if_two_chainz_orchestrated_911/,self.jokes,,He'd be called Two Planes,If Two Chainz orchestrated 9-11,0
post,3jtj08,2qh72,jokes,false,1441509964,https://old.reddit.com/r/Jokes/comments/3jtj08/yo_mama_is_so_fat/,self.jokes,,That the sorting hat put her in the waffle house!,Yo mama is so fat...,1
post,3jtil3,2qh72,jokes,false,1441509714,https://old.reddit.com/r/Jokes/comments/3jtil3/a_scotsman_is_sitting_in_a_pub/,self.jokes,,"somewhere in Scotland when an American tourist walks up to the bar. The Scotsman turns to the American, clearly drunk, and points out the window.

""Ye see that wall, right there?"" The Scotsman said in a heavy accent. ""Built that with me bare hands. But do they call me ""McGregor the Wall Builder... No...""

After another round of drinks, the Scotsman turns to the American, pointing out the window again.

""Ye see that dock there? Down by the lake?"" The Scotsman said. ""Built that with me bare hands. But do they call me 'McGregor the Dock Builder... No...""

After another round of drinks, the Scotsman turns to the American again.

""Ye fuck one sheep...""",A Scotsman is sitting in a pub...,67
post,3jtiks,2qh72,jokes,false,1441509711,https://old.reddit.com/r/Jokes/comments/3jtiks/he_was_shocked_when_this_woman_thought_hed_take/,self.jokes,,[removed],HE WAS SHOCKED WHEN THIS WOMAN THOUGHT HE’D TAKE ADVANTAGE OF HER IN A LONELY ALLEY. BUT THEN SHE SAID THIS.,0
post,3jti7h,2qh72,jokes,false,1441509504,https://old.reddit.com/r/Jokes/comments/3jti7h/what_does_the_sign_at_a_nudist_buddhist_beach_say/,self.jokes,,No [Bhikkhunis](https://en.wikipedia.org/wiki/Bhikkhuni) allowed.,What does the sign at a nudist Buddhist beach say?,14
post,3jti3p,2qh72,jokes,false,1441509451,https://old.reddit.com/r/Jokes/comments/3jti3p/a_mild_ocd_joke/,self.jokes,,"This is the joke

This is the joke


This is the joke


This is the joke


This is the joek


This is the joke



This is the joke.



This is the joke



This is the joke


This is the joke


This is the joke


This is the joke


This is the joke


This is the joke


This is the joke",A mild OCD Joke,8
post,3jthsp,2qh72,jokes,false,1441509275,https://old.reddit.com/r/Jokes/comments/3jthsp/a_bear_and_a_rabbit/,self.jokes,,"A bear and a rabbit are taking a shit in the woods. The bear turns to the rabbit and says, ""Do you have a problem with shit sticking to your fur?"" The rabbit says no.

""Great, says the bear, who then wipes his ass with the rabbit.",A bear and a rabbit,0
post,3jthhr,2qh72,jokes,false,1441509080,https://old.reddit.com/r/Jokes/comments/3jthhr/whats_it_called_when_jesus_walks_across_the_street/,self.jokes,,A cross walk,What's it called when Jesus walks across the street?,8
post,3jthe4,2qh72,jokes,false,1441509017,https://old.reddit.com/r/Jokes/comments/3jthe4/whats_the_difference_between_a_reindeer_a_knight/,self.jokes,,"The knight is slaying dragons, the reindeer is draggin' sleighs.","What's the difference between a reindeer, a knight and a cock?",0
post,3jtgy8,2qh72,jokes,false,1441508767,https://old.reddit.com/r/Jokes/comments/3jtgy8/what_did_jesus_say_after_preventing_a_crisis/,self.jokes,,[deleted],What did Jesus say after preventing a crisis?,0
post,3jtgiv,2qh72,jokes,false,1441508543,https://old.reddit.com/r/Jokes/comments/3jtgiv/my_childs_first_name/,self.jokes,,Is going to be look,My child's first name,0
post,3jtggh,2qh72,jokes,false,1441508511,https://old.reddit.com/r/Jokes/comments/3jtggh/a_group_of_philosophers_walk_into_a_bar_over/,self.jokes,,They all leave believing it's true.,"A group of philosophers walk into a bar. Over drinks, they all are trying to convince each other the statement ""All the philosophers in this group will never simultaneously believe this statement"" is false.",1
post,3jtg28,2qh72,jokes,false,1441508259,https://old.reddit.com/r/Jokes/comments/3jtg28/beethoven_was_such_a_hipster/,self.jokes,,... that he never even heard some of his own music.,Beethoven was such a hipster...,1
post,3jtfd1,2qh72,jokes,false,1441507840,https://old.reddit.com/r/Jokes/comments/3jtfd1/i_like_my_women_the_way_i_like_my_coffee/,self.jokes,,Sweet.,I like my women the way I like my coffee.,5
post,3jtf7w,2qh72,jokes,false,1441507752,https://old.reddit.com/r/Jokes/comments/3jtf7w/whats_red_but_smells_like_blue_paint/,self.jokes,,[removed],What's red but smells like blue paint?,0
post,3jtf6k,2qh72,jokes,false,1441507728,https://old.reddit.com/r/Jokes/comments/3jtf6k/reasons_why_people_want_kanye_west_as_our/,self.jokes,,"*Because people would rather have a Democratic egomaniacal maniac with no business being in politics like Kanye West, then a Republican egomaniacal maniac with no business being in politics like Donald Trump. Either I've lost faith in humanity.",Reasons Why people want Kanye West as our president over Donald Trump.,0
post,3jtei4,2qh72,jokes,false,1441507332,https://old.reddit.com/r/Jokes/comments/3jtei4/how_can_you_tell_that_your_girlfriend_is_getting/,self.jokes,,She starts fitting into your wife's clothes.,How can you tell that your girlfriend is getting fat?,2
post,3jtdy8,2qh72,jokes,false,1441506986,https://old.reddit.com/r/Jokes/comments/3jtdy8/whats_the_difference_between_jam_and_jelly/,self.jokes,,[deleted],What's the difference between Jam and Jelly?,0
post,3jtdf2,2qh72,jokes,false,1441506671,https://old.reddit.com/r/Jokes/comments/3jtdf2/i_like_my_chicken_like_i_like_my_holy_infant/,self.jokes,,"I made this up while singing silent night in the middle of field while playing capture the flag, and natural after I just ate chick tenders.",I like my chicken like I like my holy infant.. Tender and Mild,3
post,3jtcqa,2qh72,jokes,false,1441506307,https://old.reddit.com/r/Jokes/comments/3jtcqa/mr_poop/,self.jokes,,[removed],MR POOP,0
post,3jtcpt,2qh72,jokes,false,1441506299,https://old.reddit.com/r/Jokes/comments/3jtcpt/whats_the_last_thing_to_pass_through_a_gnats_mind/,self.jokes,,[deleted],What's the last thing to pass through a gnat's mind when it flies into the windshield of a car...,0
post,3jtc2u,2qh72,jokes,false,1441505915,https://old.reddit.com/r/Jokes/comments/3jtc2u/i_wish_women_had_nipples_on_their_butts/,self.jokes,,Then I could look them in the eyes as they walked away.,I wish women had nipples on their butts...,0
post,3jtbyd,2qh72,jokes,false,1441505845,https://old.reddit.com/r/Jokes/comments/3jtbyd/sister_on_her_period/,self.jokes,,"Haven't seen it on here yet, saw a similar one though.

How can you tell your sister is on her period?

Your dad's dick tastes like blood.",Sister on her period,0
post,3jtb65,2qh72,jokes,false,1441505363,https://old.reddit.com/r/Jokes/comments/3jtb65/whats_the_sin_of_unicorn_pie/,self.jokes,,[deleted],What's the sin of unicorn pie?,1
post,3jtb0i,2qh72,jokes,false,1441505259,https://old.reddit.com/r/Jokes/comments/3jtb0i/what_did_the_chef_say_when_he_was_skipped_in/,self.jokes,,Hey that's my toque!!,What did the chef say when he was skipped in rotation?,0
post,3jtafl,2qh72,jokes,false,1441504933,https://old.reddit.com/r/Jokes/comments/3jtafl/các_mẫu_đồng_hồ_nữ_đẹp_mang_đến_sự_sang_trọng_quý/,self.jokes,,đồng hồ nữ 2015,Các mẫu đồng hồ nữ đẹp mang đến sự sang trọng quý phái cho chị em,0
post,3jt9x1,2qh72,jokes,false,1441504645,https://old.reddit.com/r/Jokes/comments/3jt9x1/what_do_you_call_it_when_a_deer_knows_karate/,self.jokes,,Tae-fawn-doe,What do you call it when a deer knows karate?,6
post,3jt9vi,2qh72,jokes,false,1441504622,https://old.reddit.com/r/Jokes/comments/3jt9vi/how_many_jews_can_fit_in_a_shower/,self.jokes,,"Don't ask me, ask Hitler",How many Jews can fit in a shower?,0
post,3jt9fo,2qh72,jokes,false,1441504364,https://old.reddit.com/r/Jokes/comments/3jt9fo/how_many_cops_does_it_take_to_change_a_lightbulb/,self.jokes,,None. They just beat the room for being black.,How many cops does it take to change a lightbulb?,27
post,3jt9e4,2qh72,jokes,false,1441504339,https://old.reddit.com/r/Jokes/comments/3jt9e4/3_men/,self.jokes,,"At the National Art Gallery, in Dublin Ireland, a Canadian couple were staring at a portrait that had them completely confused.
The painting depicted three black men, totally naked, sitting on a park bench.
Two of the figures had black willies but the one in the middle had a pink one.
The curator of the gallery realized that they were having trouble interpreting the painting and offered his assessment.
He went on for over half an hour explaining how it depicted the sexual emasculation of the black man in a predominately white, patriarchal society.
“In fact,” he pointed out, “some serious critics believe that the pink also reflects the cultural and sociological oppression experienced by gay men in contemporary society.”
After the curator left, an Irish man approached the couple and said, “Would you like to know what the painting is really about?”
“Now why would you claim to be more of an expert than the curator of the gallery?” asked the husband.
“Because I’m the guy who painted it.” he replied.
”In fact, there are no black men depicted at all. They’re just three Irish coal miners. The guy in the middle went home for lunch.""
",3 Men,1
post,3jt8jc,2qh72,jokes,false,1441503879,https://old.reddit.com/r/Jokes/comments/3jt8jc/football_players_basketball_players_and_soccer/,self.jokes,,How come my girlfriend refuses to.,"Football players, basketball players and soccer players all play with balls.",0
post,3jt8fh,2qh72,jokes,false,1441503820,https://old.reddit.com/r/Jokes/comments/3jt8fh/god_will_save_me/,self.jokes,,"Heard this a while back at summer camp or something of the like. Haven't seen it on here yet.

A man is drowning in a lake. A boat drives up and the captain asks him, ""hey buddy, need any help?""  
The man responds, ""No, God will save me.""

The captain reluctantly goes about his way and a little later a speedboat drives up to the drowning man. ""Hey buddy, can I help you?""

""No, god will save me."" 

The man drowns and up in heaven he goes up to God and says, ""Hey, why didn't you save me?""

God simply replies, ""I sent you two boats, dumbass.""",God will save me,230
post,3jt89v,2qh72,jokes,false,1441503731,https://old.reddit.com/r/Jokes/comments/3jt89v/first_person_to_comment_on_this_thread_is_gau/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jt89v/first_person_to_comment_on_this_thread_is_gau/,,First person to comment on this thread is gau,20
post,3jt889,2qh72,jokes,false,1441503702,https://old.reddit.com/r/Jokes/comments/3jt889/whats_the_difference_between_chopped_beef_and_pea/,self.jokes,,"Everyone can chop beef, but no one can pee soup!",What's the difference between chopped beef and pea soup?,7
post,3jt7xa,2qh72,jokes,false,1441503544,https://old.reddit.com/r/Jokes/comments/3jt7xa/can_you_be_electrocuted_by_a_news_story/,self.jokes,,The answer may shock you. ,Can you be electrocuted by a news story?,50
post,3jt76m,2qh72,jokes,false,1441503130,https://old.reddit.com/r/Jokes/comments/3jt76m/i_cant_find_my_large_stir_fry_pan/,self.jokes,,It's like it just gets up and Woks away,I cant find my large stir fry pan,1
post,3jt72u,2qh72,jokes,false,1441503060,https://old.reddit.com/r/Jokes/comments/3jt72u/ask_someone/,self.jokes,,"If they are smart, when they inevitably say yes, ask them to spell yes. Then ask them how you would say it with an e in front of it. Enjoy as they pronounce weird words when in fact it spells eyes. ",Ask someone...,0
post,3jt6wb,2qh72,jokes,false,1441502972,https://old.reddit.com/r/Jokes/comments/3jt6wb/whats_the_average_internal_temperature_of_a/,self.jokes,,"Lukewarm, of course!",What's the average internal temperature of a Tauntaun?,2
post,3jt6k4,2qh72,jokes,false,1441502793,https://old.reddit.com/r/Jokes/comments/3jt6k4/what_did_ron_burgandy_say_when_he_dropped_his/,self.jokes,,Go fuck yourself sandy Eggo,What did Ron Burgandy say when he dropped his waffle on the beach?,13
post,3jt6ct,2qh72,jokes,false,1441502662,https://old.reddit.com/r/Jokes/comments/3jt6ct/i_painted_my_computer_black/,self.jokes,,[deleted],I painted my computer black,1
post,3jt69l,2qh72,jokes,false,1441502619,https://old.reddit.com/r/Jokes/comments/3jt69l/a_man_comes_home_to_moaning_and_groaning/,self.jokes,,"Curious, the man walks upstairs...

**Reader Reaction: UH OH! What's going to happen here? I can't imagine it being good news for the man though!**

He opens his door and he sees his wife laying there completely naked...

**Reader Reaction: Completely naked? Something fishy's going on here...**

The wife screams, ""Help! Help! I'm having a heart attack!"" In a panic, the man scrambles downstairs for the phone...

**Reader Reaction: Oh my goodness! She's having a heart att... Wait... Oh dear. I know what's going on... That's cruel for the man and a bit snide from the wife there. I hope the man finds out and kicks her into touch!""**

He sees his son and his son says, ""Hey Dad, Uncle Timmy came by earlier and he and Mom have been in the bedroom all afternoon, making weird noises."" Enraged, the man marches back upstairs...

**Reader Reaction: Hooray! Look out Uncle Timmy because here he comes! This isn't going to be pretty...""**

He marches into the room, opens the closet and sees a trembling Uncle Timmy sat there in the corner, naked. The man screams, ""My wife's having a heart attack and all you're gonna do about it is sit there butt naked in MY wardrobe?""

**Reader Reaction: Well... I wasn't expecting that! Maybe it's the best outcome, no one is hurt and everyone can move on as a family. I just hope this love affair doesn't continue!**",A man comes home to moaning and groaning,0
post,3jt523,2qh72,jokes,false,1441501969,https://old.reddit.com/r/Jokes/comments/3jt523/last_night_my_wife_said_that_our_bed_had_seen/,self.jokes,,"She's right. When she stopped at her mum's last week, I had a threesome in it on Monday and Tuesday.",Last night my wife said that our bed had seen better days.,0
post,3jt4gr,2qh72,jokes,false,1441501621,https://old.reddit.com/r/Jokes/comments/3jt4gr/who_ate_a_lot_and_conquered_rome/,self.jokes,,Atilla the Hungry.,Who ate a lot and conquered Rome?,1
post,3jt46n,2qh72,jokes,false,1441501482,https://old.reddit.com/r/Jokes/comments/3jt46n/how_did_the_stoner_die/,self.jokes,,[deleted],How did the stoner die?,0
post,3jt2n8,2qh72,jokes,false,1441500632,https://old.reddit.com/r/Jokes/comments/3jt2n8/several_days_ago_as_i_left_the_bunnings_in_rocky/,self.jokes,,[deleted],"Several days ago as I left the Bunnings in Rocky, to walk out to my ute...",2
post,3jt2jh,2qh72,jokes,false,1441500575,https://old.reddit.com/r/Jokes/comments/3jt2jh/i_like_my_women_how_i_like_my_whiskey/,self.jokes,,"12 years old and all mixed up in coke.

(sorry if its a repost, haven't seen it yet.)",I like my women how I like my whiskey.,0
post,3jt27b,2qh72,jokes,false,1441500384,https://old.reddit.com/r/Jokes/comments/3jt27b/what_do_you_call_a_mexican_baptism/,self.jokes,,Bean dip,What do you call a Mexican baptism?,2
post,3jt1a3,2qh72,jokes,false,1441499857,https://old.reddit.com/r/Jokes/comments/3jt1a3/nicki_minaj/,self.jokes,,   ,Nicki Minaj,0
post,3jt11p,2qh72,jokes,false,1441499723,https://old.reddit.com/r/Jokes/comments/3jt11p/after_being_away_from_reddit_for_a_day_how_do_you/,self.jokes,,You go to 9gag.,"After being away from Reddit for a day, how do you keep up with what you missed?",3
post,3jt0ql,2qh72,jokes,false,1441499555,https://old.reddit.com/r/Jokes/comments/3jt0ql/had_to_go_to_the_vet_so_my_dog_could_be_put_out/,self.jokes,,[deleted],Had to go to the vet so my dog could be put out of his misery...,8
post,3jt0oc,2qh72,jokes,false,1441499522,https://old.reddit.com/r/Jokes/comments/3jt0oc/a_man_on_a_plane/,self.jokes,,"A man boarded an airplane and took his seat. As he settled in, he glanced Up and saw the most beautiful woman boarding the plane. He soon realized She was heading straight towards his seat. As fate would have it, she took The seat right beside his. Eager to strike up a conversation he blurted out, “Business trip or pleasure?”
She turned, smiled and said, “Business. I’m going to the Annual Nymphomaniacs of America Convention in Boston.""
He swallowed hard. Here was the most gorgeous woman he had ever seen Sitting next to him, and she was going to a meeting of nymphomaniacs!
Struggling to maintain his composure, he calmly asked, “What’s your Business at this convention?”
“Lecturer,” she responded. “I use information that I have learned from my Personal experiences to debunk some of the popular myths about sexuality.”
“Really?” he said. “And what kind of myths are there?”
“Well,” she explained, “one popular myth is that African-American men are The most well-endowed of all men, when in fact it is the Native American Indian who is most likely to possess that trait. Another popular myth is That Frenchmen are the best lovers, when actually it is men of Mexican Descent who are the best. I have also discovered that the lover with Absolutely the best stamina is the Southern Redneck.”
Suddenly the woman became a little uncomfortable and blushed.. “I’m Sorry,” she said, “I shouldn't really be discussing all of this with you. I don’t Even know your name.”
“Tonto,” the man said, “Tonto Gonzales, but my friends call me Bubba"".",A man on a plane,261
post,3jt0fq,2qh72,jokes,false,1441499393,https://old.reddit.com/r/Jokes/comments/3jt0fq/there_were_these_two_guys_in_a_lunatic_asylum/,self.jokes,,"See, there were these two guys in a lunatic asylum...and one night, one night they decide they don't like living in an asylum any more. They decide they're going to escape! So, like, they get up onto the roof and there, just across this narrow gap, they see the rooftops of the town, stretching away in the moonlight...stretching away to freedom. Now, the first guy, he jumps right across with no problem. But his friend, his friend daren't make the leap. Y'see...y'see, he's afraid of falling. So then, the first guy has an idea...He says 'Hey! I have my flashlight with me! I'll shine it across the gap between the buildings. You can walk along the beam and join me!' B-but the second guy just shakes his head. He suh-says... he says 'What do you think I am? Crazy? You'd turn it off when I was half way across!'
Then the Batman stopped them. ",There were these two guys in a lunatic asylum,0
post,3jt0ff,2qh72,jokes,false,1441499389,https://old.reddit.com/r/Jokes/comments/3jt0ff/what_is_the_bird_synonymous_with_abstinence/,self.jokes,,The Swallow,What is the bird synonymous with abstinence,1
post,3jt011,2qh72,jokes,false,1441499190,https://old.reddit.com/r/Jokes/comments/3jt011/why_did_the_plane_crash_into_the_mountain/,self.jokes,,Because the pilot was a loaf of bread. ,Why did the plane crash into the mountain?,0
post,3jszl1,2qh72,jokes,false,1441498954,https://old.reddit.com/r/Jokes/comments/3jszl1/life_is_like_a_box_of_chocolates/,self.jokes,,neither lasts long for a fat person,Life is like a box of chocolates,140
post,3jszhz,2qh72,jokes,false,1441498910,https://old.reddit.com/r/Jokes/comments/3jszhz/what_did_the_locomotive_conductor_crave_once_he/,self.jokes,,traaaiins...,what did the locomotive conductor crave once he became a zombie?,2
post,3jsz6j,2qh72,jokes,false,1441498720,https://old.reddit.com/r/Jokes/comments/3jsz6j/i_came_home_from_work_early_today_and_caught_my/,self.jokes,,"""That's disgusting"" I said, ""I'm meant to be eating that tonight, now it's going to taste like salad.""",I came home from work early today and caught my daughter masturbating with a cucumber,0
post,3jsxjg,2qh72,jokes,false,1441497791,https://old.reddit.com/r/Jokes/comments/3jsxjg/an_old_man_and_a_teenager_are_talking_in_the/,self.jokes,,"The old man says, ""It's your generation that's destroying our society.""

**Reader Reaction: Ugh! That nasty cynical old man! That's obviously not true! I hope he gets his comeuppance!**

The teenager replies, ""Man, if I had a dollar for every time someone said that to me, I'd have enough money to buy a house in the economy YOU destroyed!""

**Reader Reaction: OOOH! Take that you uncouth old man! I'm glad he got found out and we all learned a valuable lesson today that nobody is perfect!**",An old man and a teenager are talking in the street,0
post,3jsxew,2qh72,jokes,false,1441497728,https://old.reddit.com/r/Jokes/comments/3jsxew/i_didnt_really_want_to_go_to_the_seafood_buffet/,self.jokes,,...but I just went for the halibut,I didn't really want to go to the seafood buffet...,24
post,3jswgw,2qh72,jokes,false,1441497208,https://old.reddit.com/r/Jokes/comments/3jswgw/a_man_is_walking_home_from_the_market_with_three/,self.jokes,,"Fumbling with everything, he asks a lady on the street to please hold one of the pigs for him while he figures out how to carry it all.


""No! You could *rape* me!""


""Lady, how in the world could I rape you holding two pigs and a wash tub?""


Lady thinks a minute and says, ""Well, you could put one under the wash tub, make me stand on top of it, you hold one and I could hold the other.""



(Thanks, Dad. RIP in peace.)",A man is walking home from the market with three pigs and a wash tub.,7
post,3jswe2,2qh72,jokes,false,1441497165,https://old.reddit.com/r/Jokes/comments/3jswe2/whats_the_difference_between_a_garbanzo_bean_and/,self.jokes,,I never had a garbanzo bean on my face.,What's the difference between a garbanzo bean and a chick pea?,17
post,3jswas,2qh72,jokes,false,1441497116,https://old.reddit.com/r/Jokes/comments/3jswas/what_happens_when_you_throw_a_piano_down_a_mine/,self.jokes,,A flat miner.,What happens when you throw a piano down a mine shaft?,2
post,3jsw0j,2qh72,jokes,false,1441496964,https://old.reddit.com/r/Jokes/comments/3jsw0j/what_do_you_call_a_black_person/,self.jokes,,[removed],what do you call a black person?,1
post,3jsvt1,2qh72,jokes,false,1441496839,https://old.reddit.com/r/Jokes/comments/3jsvt1/there_is_a_monkey_in_a_bar_a_sign_says_feel_free/,self.jokes,,"A man sees the sign and decides to feed the monkey a peanut. He gives the peanut to the monkey.

The monkey shoves the peanut up it's ass, then takes the peanut out and eats it.

Amused, the man asks the bartender:"" Dude, why does that monkey do that?""

The bartender laughs:"" He's been like that ever since he ate the cue ball.""","There is a monkey in a bar. A sign says ""feel free to feed the monkey.""",7
post,3jsvre,2qh72,jokes,false,1441496812,https://old.reddit.com/r/Jokes/comments/3jsvre/what_do_you_say_to_guy_who_is_wearing_an_apple/,self.jokes,,[deleted],What do you say to guy who is wearing an apple watch?,1
post,3jsvfl,2qh72,jokes,false,1441496628,https://old.reddit.com/r/Jokes/comments/3jsvfl/whats_green_and_has_wheels/,self.jokes,,[deleted],What's green and has wheels?,0
post,3jsuul,2qh72,jokes,false,1441496336,https://old.reddit.com/r/Jokes/comments/3jsuul/livewisconsin_vs_alabama_live_stream_ncaa_college/,self.jokes,,[removed],LIVE]]@.Wisconsin vs Alabama Live Stream.. NCAA.. College.. Football.. Alabama vs Wisconsin Streaming..Sept..5th..,1
post,3jsunr,2qh72,jokes,false,1441496241,https://old.reddit.com/r/Jokes/comments/3jsunr/an_old_man_and_a_teenager_are_talking_on_the/,self.jokes,,[removed],An old man and a teenager are talking on the street (INCLUDES READER REACTION FEATURE),1
post,3jsui5,2qh72,jokes,false,1441496160,https://old.reddit.com/r/Jokes/comments/3jsui5/what_does_op_and_digiorno_have_in_common/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jsui5/what_does_op_and_digiorno_have_in_common/,,What does OP and DiGiorno have in common?,54
post,3jsu9m,2qh72,jokes,false,1441496037,https://old.reddit.com/r/Jokes/comments/3jsu9m/what_happens_if_you_run_out_of_prisoners_at/,self.jokes,,[deleted],What happens if you run out of prisoners at Guantanamo Bay?,2
post,3jstt5,2qh72,jokes,false,1441495822,https://old.reddit.com/r/Jokes/comments/3jstt5/the_one_thing_that_i_excel_at/,self.jokes,,is spreadsheets. ,The one thing that I excel at...,2
post,3jstrh,2qh72,jokes,false,1441495801,https://old.reddit.com/r/Jokes/comments/3jstrh/parking_spot/,self.jokes,,"An old man was driving downtown in his Bentley. He drove around for 45 minutes until he saw a spot on the side of the street. As the spot freed up another man in a Lamborghini slides in and takes it before the old man can. As the other drive stepped out of his vehicle, he looks at the old man and says: ""You need to be fast to do that!"". The old man takes a second and slams his Bentley into the Lambo, pushing it out of the spot. he then backs in and with a wrecked front end. With calm composure he steps out of his car and looks at the Lambo driver and says: ""You need to be rich to do that!"" and walks away.",Parking spot,1
post,3jst0v,2qh72,jokes,false,1441495412,https://old.reddit.com/r/Jokes/comments/3jst0v/what_porn_do_vampires_love/,self.jokes,,Fangbang,What porn do vampires love?,2
post,3jssx0,2qh72,jokes,false,1441495356,https://old.reddit.com/r/Jokes/comments/3jssx0/a_young_man_has_sex_for_the_first_time/,self.jokes,,"The young man was very nervous about having sex with his girlfriend for the very first time, because he was convinced that his penis would be too small.

Eventually he realized that he could not postpone it forever and he nervously invited her over to his house.

Hesitatingly he started to take off his clothes and after that he dimmed the lights. Very carefully he started taking off her clothes and he started stroking her. 

Finally he nervously nestled his erection inside her hand, hoping she didn't realize how small it was.

""No thank you,"" she said, ""I don't smoke.""",A young man has sex for the first time,3829
post,3jsrg6,2qh72,jokes,false,1441494587,https://old.reddit.com/r/Jokes/comments/3jsrg6/husband_and_wife_were_watching_national_geographic/,self.jokes,,[removed],Husband and wife were watching National Geographic,0
post,3jsqnm,2qh72,jokes,false,1441494189,https://old.reddit.com/r/Jokes/comments/3jsqnm/i_finally_got_around_to_reading_that_book_on/,self.jokes,,It's about time.,I finally got around to reading that book on watches I got last year,4
post,3jsqg1,2qh72,jokes,false,1441494084,https://old.reddit.com/r/Jokes/comments/3jsqg1/a_woman_is_complaining_to_her_neighbor/,self.jokes,,"A woman is complaining to her neighbor:
- My husband is 300% impotent.
- A few days ago you told me 100%, not 300%.
- Well, yesterday he fell down the stairs, broke his finger and bit his tongue.",A woman is complaining to her neighbor,14
post,3jsq4q,2qh72,jokes,false,1441493932,https://old.reddit.com/r/Jokes/comments/3jsq4q/whats_the_popes_least_favorite_human_bone/,self.jokes,,The blasphemur.,What's the Pope's least favorite human bone?,0
post,3jspsb,2qh72,jokes,false,1441493744,https://old.reddit.com/r/Jokes/comments/3jspsb/you_hear_about_the_chinese_godfather/,self,self,,You hear about the Chinese godfather?,1
post,3jspjn,2qh72,jokes,false,1441493607,https://old.reddit.com/r/Jokes/comments/3jspjn/how_do_you_find_a_blind_man_in_a_nudist_colony/,self.jokes,,Its not hard.,How do you find a blind man in a nudist colony?,2
post,3jsp3i,2qh72,jokes,false,1441493384,https://old.reddit.com/r/Jokes/comments/3jsp3i/a_man_went_to_a_farm_after_being_lost/,self.jokes,,"Once he arrive to the door he knocked 3 times exactly . 

No answer , so he knocked 3 more times . 

Still no answer , the man was getting furious so he decided to kick the door instead , by his suprise an old man answered 

The old man then aproached him and said ""yes sir , sorry I don't have my hearing aid I hope you didn't wait too long""

He then proceeds to invite him in for supper , the old man sat down and so did he . While he was eating away , old man starts asking questions . 

""So where are you from boy"" 

""Oh I don't really wanna talk about that""

""well can you atleast tell me why you are here"" the old man said 

Quickly the young one said ""I was lost for 2 days , I needed food and water "" 

The old man laughing , wondering how he got lost in these woods then says ""what's your name young one ?""

The young boy replies ""JOOOOOOOOOOHN CENAAAAAAAAAAAA""

DOOOOT DOOT DOOT DOOT

Edit : sorry I'm tired,  don't kill me",A man went to a farm after being lost,0
post,3jsooa,2qh72,jokes,false,1441493163,https://old.reddit.com/r/Jokes/comments/3jsooa/dark_humor_is_like_food/,self.jokes,,Not everyone gets it.,Dark humor is like food.,20
post,3jso96,2qh72,jokes,false,1441492958,https://old.reddit.com/r/Jokes/comments/3jso96/i_bought_my_shoes_from_a_drug_dealer/,self.jokes,,"I don't know what he laced them with, but I've been trippin' all day. ",I bought my shoes from a drug dealer.,23
post,3jso81,2qh72,jokes,false,1441492940,https://old.reddit.com/r/Jokes/comments/3jso81/for_my_cake_day_i_present_to_you_one_of_my/,self.jokes,,[deleted],For my cake day I present to you one of my favorites - What type of gas do you fart?,0
post,3jsn07,2qh72,jokes,false,1441492351,https://old.reddit.com/r/Jokes/comments/3jsn07/i_saw_a_bloke_let_his_dog_walk_straight_out_in/,self.jokes,,"The cruel cunt didn't even flinch when it was killed. He was too busy standing round, trying to look cool in his sunglasses, swinging his walking stick about like he didn't care.",I saw a bloke let his dog walk straight out in front of a lorry this morning.,0
post,3jslb8,2qh72,jokes,false,1441491542,https://old.reddit.com/r/Jokes/comments/3jslb8/what_do_you_call_a_blind_alien/,self.jokes,,[deleted],What do you call a blind alien?,1
post,3jsl31,2qh72,jokes,false,1441491432,https://old.reddit.com/r/Jokes/comments/3jsl31/do_you_know_why_one_side_of_the_v_is_slightly/,self.jokes,,Because there are more birds on that side.,Do you know why one side of the V Is slightly larger when birds fly together?,3
post,3jskop,2qh72,jokes,false,1441491249,https://old.reddit.com/r/Jokes/comments/3jskop/whats_the_difference_between_a_cheese/,self.jokes,,[deleted],What's the difference between a cheese?,0
post,3jskdn,2qh72,jokes,false,1441491115,https://old.reddit.com/r/Jokes/comments/3jskdn/what_cheese_do_you_take_with_you_on_a_bear_hunt/,self.jokes,,Camembert.,What cheese do you take with you on a bear hunt?,0
post,3jsk4e,2qh72,jokes,false,1441490993,https://old.reddit.com/r/Jokes/comments/3jsk4e/little_johnny/,self.jokes,,"Little Johnny says to the teacher..

Miss, Miss I need to do a piss! The teacher says ' Johnny, the proper term is urinate. I want you to go to the toilet and when you come back i want you to use urinate in a sentence.'

Little Johnny goes to the toilet and rushes back. Teacher: ok Johnny, use urinate in a sentence. Johnny flashes back, ""ok miss, urinate, but if you had bigger tits, you'd be a 10!""",Little Johnny...,110
post,3jsjti,2qh72,jokes,false,1441490841,https://old.reddit.com/r/Jokes/comments/3jsjti/dad_jokes_for_fathers_day/,self.jokes,,"As its Father's Day (in Australia at least), here's a thread for all our favourite Dad Jokes

How many tickles does it take to make an octopus laugh? Ten tickles


Happy Dad Joke Day!",Dad jokes for Father's Day,9
post,3jsj3n,2qh72,jokes,false,1441490496,https://old.reddit.com/r/Jokes/comments/3jsj3n/freedom_units_are_measured_in/,self.jokes,,Caliber.,Freedom Units are Measured In...,2
post,3jsi9m,2qh72,jokes,false,1441490128,https://old.reddit.com/r/Jokes/comments/3jsi9m/what_did_the_pirate_say_when_he_turned_80/,self.jokes,,Aye matey,What did the pirate say when he turned 80?,1
post,3jsh2q,2qh72,jokes,false,1441489576,https://old.reddit.com/r/Jokes/comments/3jsh2q/a_mum_and_dad_is_sitting_at_the_table_with_their/,self.jokes,,[deleted],A mum and dad is sitting at the table with their blind son discussing a relevant political situation.,2
post,3jsgre,2qh72,jokes,false,1441489428,https://old.reddit.com/r/Jokes/comments/3jsgre/teacher_translate_this_russian_sentence_into/,self.jokes,,"Teacher Translate This Russian Sentence into English
Она приезжает сюда слепой ( She is coming here )
Russian Student. A blind Girl is Sleeping here",Teacher Translate This Russian Sentence into English,0
post,3jsgqa,2qh72,jokes,false,1441489411,https://old.reddit.com/r/Jokes/comments/3jsgqa/what_do_you_call_a_chinese_man_sitting_on_a_wall/,self.jokes,,Ray ling,What do you call a Chinese man sitting on a wall?,0
post,3jsfyz,2qh72,jokes,false,1441489051,https://old.reddit.com/r/Jokes/comments/3jsfyz/in_the_jungle_the_mighty_jungle_the_lions/,self.jokes,,"A male and female lion are taking a siesta I'm the hot savanna heat when a jackal appear.
He walks back and forth and look at the female lion and start to curse: ho, cunt, bitch. 
Furious, she stands on all four ready to leap when the male lion says, don't do it.
She puts a paw forward and the jackal runs away.
She lies down and before you know it the jackal is back.
Cunt, slut, ho...
Once again she stands up and the other lion goes,
Don't do it, trust me.
The jackal just keep shooting off his foul mouth and she just snaps and starts to chase the little fucker.
After a minute of running the jackal runs inside a small drainage pipe and the lioness follows and gets stuck.
The jackal comes out from the other side, circles around and comes up behind her, lifts up her tail and does his business... 
After a couple of hours she comes back, limping and groggy.
The male lion looks at her and says, he took you to the pipe ehhh.","In the jungle, the mighty jungle, the lions...",4
post,3jsfe4,2qh72,jokes,false,1441488790,https://old.reddit.com/r/Jokes/comments/3jsfe4/whats_an_owls_favorite_subject/,self.jokes,,Owlgebra,What's an owl's favorite subject?,3
post,3jsf7h,2qh72,jokes,false,1441488707,https://old.reddit.com/r/Jokes/comments/3jsf7h/what_do_you_get_when_you_mix_a_dog_and_a_tulip/,self.jokes,,A collieflower ,What do you get when you mix a dog and a tulip?,1
post,3jseuj,2qh72,jokes,false,1441488543,https://old.reddit.com/r/Jokes/comments/3jseuj/whats_a_caterpillar_afraid_of/,self.jokes,,"A dogerpillar


(Thank you Laffy Taffy for the ~~worst~~ best joke I've ever heard)",What's a caterpillar afraid of?,0
post,3jseo2,2qh72,jokes,false,1441488458,https://old.reddit.com/r/Jokes/comments/3jseo2/two_guys_in_an_asylum_decide_one_night_theyre/,self.jokes,,"However, the first guy has an idea...
He says ""Hey! I got my flashlight! I'll shine it across the gap between the buildings. You can walk along the beam and join me!"" 

The second guy just shakes his head and says: ""Wh-what do you think I am? Crazy? You'd turn off the light when I was halfway across!"" ","Two guys in an asylum decide one night they're sick of living there, and decide to escape. They make their way to the roof, and just across this tiny gap are the rooftops of the town, glowing in the moon light. Freedom The first guy jumps right across but his pal didn't dare for fear of falling.",6
post,3jse73,2qh72,jokes,false,1441488255,https://old.reddit.com/r/Jokes/comments/3jse73/the_day_after_his_wife_disappeared_in_a_kayaking/,self.jokes,,"...An Anchorage man answered his door to find two grim-faced Alaska State Troopers.
""We're sorry, Mr. Wilkens, but we have some information about your wife,"" said one trooper.
""Tell me! Did you find her?!"" Wilkens shouted.
The troopers looked at each other, One said, ""We have some bad news, some good news, and some really great news. Which do you want to hear first?""
Fearing the worst, an ashen Mr. Wilkens said, ""Give me the bad news first.""
The trooper said, ""I'm sorry to tell you, sir, but this morning we found your wife's body in Kachemak Bay.""
""Oh, no!"" exclaimed Wilkens. Swallowing hard, he asked, ""What's the good news?""
The trooper continued, ""When we pulled her up, she had 12 twenty-five pound king crabs and 6 good-sized Dungeness crabs clinging to her.""
Stunned, Mr. Wilkens demanded, ""If that's the good news, what's the great news?""
The trooper said, ""Tomorrow, we're going to pull her up again!""",The day after his wife disappeared in a kayaking accident....,58
post,3jsdfl,2qh72,jokes,false,1441487925,https://old.reddit.com/r/Jokes/comments/3jsdfl/why_will_you_never_starve_in_the_desert/,self.jokes,,[deleted],Why will you never starve in the desert?,1
post,3jsc3n,2qh72,jokes,false,1441487328,https://old.reddit.com/r/Jokes/comments/3jsc3n/i_told_my_friend_to_not_worry_about_being_hungry/,self.jokes,,Because of all the sand which is there.,I told my friend to not worry about being hungry at the beach.,23
post,3jsbm4,2qh72,jokes,false,1441487088,https://old.reddit.com/r/Jokes/comments/3jsbm4/what_pick_up_line_does_jared_from_subway_use/,self.jokes,,[deleted],What pick up line does Jared from Subway use?,0
post,3jsbjb,2qh72,jokes,false,1441487051,https://old.reddit.com/r/Jokes/comments/3jsbjb/what_do_you_call_a_reptile_that_loves_putting/,self.jokes,,a segreGATOR,What do you call a reptile that loves putting things in groups?,2
post,3jsbhj,2qh72,jokes,false,1441487032,https://old.reddit.com/r/Jokes/comments/3jsbhj/on_leftovers/,self.jokes,,[removed],On Leftovers,1
post,3jsak0,2qh72,jokes,false,1441486610,https://old.reddit.com/r/Jokes/comments/3jsak0/i_never_understood_why_people_associate_sign/,self.jokes,,[deleted],I never understood why people associate sign language with deaf people,0
post,3jsaee,2qh72,jokes,false,1441486541,https://old.reddit.com/r/Jokes/comments/3jsaee/enjoy_southern_illinois_vs_indiana_live_hd_tv/,self.jokes,,[removed],Enjoy Southern Illinois vs Indiana live HD TV NCAA Footba...,1
post,3jsa7k,2qh72,jokes,false,1441486447,https://old.reddit.com/r/Jokes/comments/3jsa7k/a_really_funny_joke_i_thought_about_link_is_in/,self.jokes,,[Hope you like it!](http://zelda.wikia.com/wiki/Link),"A really funny joke I thought about, link is in the description.",1
post,3js9pv,2qh72,jokes,false,1441486209,https://old.reddit.com/r/Jokes/comments/3js9pv/how_to_get_republicans_to_be_cool_with_gay/,self.jokes,,[deleted],How to get Republicans to be cool with Gay Marriage in America,0
post,3js9mm,2qh72,jokes,false,1441486163,https://old.reddit.com/r/Jokes/comments/3js9mm/how_do_you_eat_a_computer/,self.jokes,,byte by byte. ,How do you eat a computer?,20
post,3js9mi,2qh72,jokes,false,1441486161,https://old.reddit.com/r/Jokes/comments/3js9mi/a_man_going_through_a_divorce/,self.jokes,,"A man going through a divorce....Is walking on the beach. He comes across something in the sand.It's a lamp! The man rubs it and a genie appears!""I am so and so(insert name)!"", said the genie. ""I can grant you three wishes of whatever worldly possession imaginable, BUT since you rubbed my lamp. I now have a bond with you that allows me to see your life and try to fulfill whatever your heart desires.."" ""That being said, your soon to be ex wife will receive double what you wish for! I know it seems unfair, but rules are rules."" The man begins to thinks very intensely. Then jumps up, "" I know!""""For my first wish, I wish for 10 million dollars"", said the man.""Remember"", said the genie. ""Your wife gets double!"" The man nods in agreement. POOF! Now the man has 10 million dollars in the bank.""Now your second wish!""demanded the genie.""I wish for a mansion by the ocean!""POOF! They appear in a beautiful mansion!""Now....Tell me what your last wish is..."", said the genie..""I wish to be beaten half to death!!""TR;DR Find a lamp with a genie in it? Choose your wishes wisely...",A man going through a divorce...,1
post,3js8yw,2qh72,jokes,false,1441485850,https://old.reddit.com/r/Jokes/comments/3js8yw/2_lepers_playing_poker/,self.jokes,,"1 throws his hand in, the other laughs his head off. ",2 lepers playing poker...,4
post,3js8kg,2qh72,jokes,false,1441485649,https://old.reddit.com/r/Jokes/comments/3js8kg/two_guys_are_walking_down_the_street_when_a/,self.jokes,," Just then one guy turns to the other and hands him a bill. “Here’s that $20 I owe you,” he says.",Two guys are walking down the street when a mugger approaches them and demands their money. They both grudgingly pull out their wallets and begin taking out their cash..,4
post,3js7ro,2qh72,jokes,false,1441485269,https://old.reddit.com/r/Jokes/comments/3js7ro/how_do_you_punish_a_rock/,self.jokes,,[deleted],How do you punish a rock?,4
post,3js7dq,2qh72,jokes,false,1441485085,https://old.reddit.com/r/Jokes/comments/3js7dq/the_best_part_of_swiss_cheese/,self.jokes,,Is the holes,The best part of Swiss cheese,0
post,3js784,2qh72,jokes,false,1441485009,https://old.reddit.com/r/Jokes/comments/3js784/why_was_six_afraid_of_seven/,self.jokes,,"Because it saw seven set a hobo on fire and masturbate on his charred corpse.

(Source: Patton Oswalt)",Why was six afraid of seven?,7
post,3js70j,2qh72,jokes,false,1441484917,https://old.reddit.com/r/Jokes/comments/3js70j/why_is_no_one_friends_with_dracula/,self.jokes,,Cause hes a pain in the neck.,Why is no one friends with Dracula?,7
post,3js6hm,2qh72,jokes,false,1441484683,https://old.reddit.com/r/Jokes/comments/3js6hm/why_do_most_newfie_men_have_beards_or_mustaches/,self.jokes,,They wanna look just like their mothers.,Why do most newfie men have beards or mustaches?,2
post,3js67h,2qh72,jokes,false,1441484556,https://old.reddit.com/r/Jokes/comments/3js67h/what_do_you_call_the_dapper_bouncer_at_a_coin_op/,self.jokes,,"The Deter Gent.

;D",What do you call the dapper bouncer at a coin op laundromat?,1
post,3js63l,2qh72,jokes,false,1441484503,https://old.reddit.com/r/Jokes/comments/3js63l/whats_the_difference_between_a_black_man_and_an/,self.jokes,,One is a nerdy digger.,What's the difference between a black man and an archealogist?,4
post,3js57t,2qh72,jokes,false,1441484116,https://old.reddit.com/r/Jokes/comments/3js57t/ed_the_rancher_drives_to_buy_a_new_tractor_and/,self.jokes,,"Very nervous, he goes along to the lingerie shop and walks up to the pretty salesgirl.

”Can I help you, sir?” asks the girl.

Ed points to a bra on a dummy, blushes, and stammers, ”I wanna buy one of those things.”

”Certainly, sir,” replies the girl. ”What size?”

”Size?” gasps Ed. ”Ah! My God! I don’t know!”

”Well,” says the girl, helpfully, ”are they like coconuts?”

”Oh no!” replies Ed.

”Well then, are they like grapefruits?” she asks.

”No, not at all,” replies Ed.

”Oranges then,” suggests the girl.

”No,” replies Ed.

”Lemons?” she asks.

”Lemons?” repeats Ed. ”Ah, no!”

”Well then, how about eggs,” suggests the girl.

”Eggs... yes, eggs!” says Ed, confidently – ”fried eggs!”","Ed, the rancher, drives to buy a new tractor, and wants to get a present for Mabel, his wife.",0
post,3js516,2qh72,jokes,false,1441484035,https://old.reddit.com/r/Jokes/comments/3js516/whats_the_difference_between_a_dirty_bus_stop_and/,self.jokes,,"one's a crusty bus station, and the other's a busty crustacean.",Whats the difference between a dirty bus stop and a lobster with breast implants?,18
post,3js4qq,2qh72,jokes,false,1441483902,https://old.reddit.com/r/Jokes/comments/3js4qq/come_on_guys_give_us_your_best_your_momma_jokes/,self.jokes,,"* Your momma is so fat that NASA uses her for gravity assist maneuvers.
* Your momma is so fat that her belly button is an event horizon.
* Your momma is so fat and old that once when she tripped and fell over , the moon was created.
* Your momma is so fat that I can see what's behind her due to gravitational lensing.
* Your momma is so fat that she is considered to be a viable candidate for the recolonization of the human race once we have depleted our planet of it's natural resources.
* Your momma is so fat that she doesn't go to the beach, the beach comes to her.
* Your momma is so fat that when aliens tried to abduct her, their tractor beam broke down.","Come on guys! Give us your best ""Your Momma"" jokes!",0
post,3js3u2,2qh72,jokes,false,1441483528,https://old.reddit.com/r/Jokes/comments/3js3u2/if_memes_were_horses/,self.jokes,,"4chan would give birth to it.

Reddit would kill it.

9Gag would hump its dead body.

Facebook would dig up its corpse and attempt to turn its remains into Frankenstein.",If Memes Were Horses,2
post,3js3sb,2qh72,jokes,false,1441483510,https://old.reddit.com/r/Jokes/comments/3js3sb/president_kanye_west/,self.jokes,,[deleted],President Kanye West.,0
post,3js3qo,2qh72,jokes,false,1441483493,https://old.reddit.com/r/Jokes/comments/3js3qo/what_do_you_call_a_conservative_acting_as_a_mole/,self.jokes,,A decepti-con.,What do you call a conservative acting as a mole in the Democratic party?,2
post,3js3ks,2qh72,jokes,false,1441483424,https://old.reddit.com/r/Jokes/comments/3js3ks/surfs_up/,self.jokes,,"A Californian surfer visiting Australia was having a good time catching the breakers at resorts along the Gold Coast, but wanted a special experience. He wanted to surf a beach where nobody, or almost nobody, goes.

So he gets in the car, drives north. At the first remote beach he hits, he has his board in hand as he's walking toward the water, when one of the locals warns him: ""you don't want to be surfing here, mate: there's too many sharks"".

So he heeds the warning, and drives to one remote beach after another - and it's always the same warning: there's too many sharks.

Finally, he finds a perfect beach. It's so perfect, film editors would cut it out because the audience would never believe it's real. He asks the first person he meets if there are any sharks here, and was told, no.

Two more locals give him the same answer: no sharks here. So he splashes into the water and paddles out toward the breakers, when the alarm goes off in his head. This is a perfect beach, the water temperature's perfect, the breakers are to die for... and not only are there no surfers, nobody is in the water. Something's got to be wrong.

So he turns his head and cries out to a sunbather catching a tan: ""Hey, why aren't there any sharks at this beach?""

And the guy answers: ""because they're bloody afraid of the crocodiles, mate!""",Surf's up?,5
post,3js35j,2qh72,jokes,false,1441483246,https://old.reddit.com/r/Jokes/comments/3js35j/how_do_you_approach_an_angry_welsh_cheese/,self.jokes,,Caerphilly.,How do you approach an angry Welsh cheese?,3
post,3js2m4,2qh72,jokes,false,1441483029,https://old.reddit.com/r/Jokes/comments/3js2m4/what_do_you_call_a_cross_between_a_joke_and_a/,self.jokes,,[deleted],What do you call a cross between a joke and a rhetorical question?,0
post,3js272,2qh72,jokes,false,1441482848,https://old.reddit.com/r/Jokes/comments/3js272/your_mommas_so_fat_they_use_her_as_the_wrecking/,self.jokes,,[deleted],Your momma's so fat they use her as the wrecking ball.,0
post,3js1hw,2qh72,jokes,false,1441482530,https://old.reddit.com/r/Jokes/comments/3js1hw/a_drunk_walk_into_a_saloon/,self.jokes,,"With no money in his pockets he start to beg.
With no luck he begins to get desperate and yells out ""I’ll do anything"".
The bartender looks at him and says:
If you take a sip from the spitoon then I’ll give you a bottle.
The desperate man walked back and forth a couple of times before he decided to do it, he walked up to the spitoon, lifted it up and started to drink, one chug after another until it was empty.
The bartender looks at him, gives him the bottle and asks:
Why did you drink it all up? I said a sip was enough.
The drunk looked back at him and said:
I was planning to but the pieces of mucus just would not separate.",A drunk walk into a saloon!,2
post,3js1cl,2qh72,jokes,false,1441482463,https://old.reddit.com/r/Jokes/comments/3js1cl/little_johnny_with_teacher/,self.jokes,,"Little Johnny: Teacher, can I go to the bathroom? 
Teacher: Little Johnny, MAY I go to the bathroom? 
Little Johnny: But I asked first",Little Johnny With Teacher,1
post,3js17j,2qh72,jokes,false,1441482401,https://old.reddit.com/r/Jokes/comments/3js17j/why_is_germany_taking_in_immigrants/,self.jokes,,because they have the camps.,Why is Germany taking in immigrants,0
post,3js101,2qh72,jokes,false,1441482296,https://old.reddit.com/r/Jokes/comments/3js101/whats_do_a_baby_and_old_people_have_in_common/,self.jokes,,They both get ditched in the park,Whats do a baby and old people have in common?,0
post,3js0dw,2qh72,jokes,false,1441482000,https://old.reddit.com/r/Jokes/comments/3js0dw/whats_better_than_roses_on_your_piano/,self.jokes,,Tulips on your organ.,What's better than roses on your piano?,3
post,3jrza5,2qh72,jokes,false,1441481463,https://old.reddit.com/r/Jokes/comments/3jrza5/a_woman_is_in_bed_with_her_lover_who_also_happens/,self.jokes,,"They had sex for hours, and afterwards, while they're just laying there, the phone rings.
Since it is the woman's house, she picks up the receiver. Her lover looks over at her and listens, only hearing her side of the conversation... She is speaking in a cheery voice) ""Hello? Oh, hi. I'm... so glad that you called. Really? That's wonderful. I am so happy for you. That sounds terrific. Great! Thanks. Okay. Bye.""
She hangs up the telephone and her lover asks, ""Who was that?""
""Oh"" she replies, ""that was my husband telling me all about the wonderful time he's having on his fishing trip with you.""",A woman is in bed with her lover who also happens to be her husband's best friend.,43
post,3jrz9m,2qh72,jokes,false,1441481455,https://old.reddit.com/r/Jokes/comments/3jrz9m/two_hobos_walking_along_the_tracks/,self.jokes,,"One hobo turns to the other and asks: ""You stink! Did you shit your pants? ""

The other hobo says emphatically: ""No! ""

An hour later as the day gets hotter the first hobo says: "" You STILL stink, and it's *worse*! Tell me the truth. . DID YOU SHIT YOUR PANTS?!""

The second hobo once again denies it. 

Finally,  as the day's heat reaches is peak and the smell becomes overwhelming, the first hobo just reaches over and yanks the other hobos pants down where he sees his underwear is packed with so much shit, it's oozing from the seams. The first hobo says: ""I can SEE the shit in your pants!  Why did you say you didn't shit your pants?!?""

The second hobo says: ""I thought you meant *today*!""",Two hobos walking along the tracks.....,2
post,3jryb8,2qh72,jokes,false,1441480974,https://old.reddit.com/r/Jokes/comments/3jryb8/knock_knock/,self.jokes,,"Who's there?

Banana

Banana who?

KEVIN!",Knock knock.,0
post,3jrwt3,2qh72,jokes,false,1441480319,https://old.reddit.com/r/Jokes/comments/3jrwt3/whats_the_difference_between_a_high_school_girls/,self.jokes,,Pigmies are a cunning bunch of runts. ,What's the difference between a High School girls track team and a tribe of pigmy?,5
post,3jrwdm,2qh72,jokes,false,1441480148,https://old.reddit.com/r/Jokes/comments/3jrwdm/some_aquatics_mammals_escaped_from_the_zoo_the/,self.jokes,,it was otter chaos.,Some aquatics mammals escaped from the zoo the other day..,1
post,3jrvuo,2qh72,jokes,false,1441479912,https://old.reddit.com/r/Jokes/comments/3jrvuo/how_can_you_tell_the_difference_between_a/,self.jokes,,"One you'll see in a while, the other you'll see later.
Credit to Mitch hedburg",How can you tell the difference between a crocodile and an alligator?,9
post,3jrvi3,2qh72,jokes,false,1441479762,https://old.reddit.com/r/Jokes/comments/3jrvi3/my_spanish_teacher_asked_me_to_turn_in_my_essay/,self.jokes,,[deleted],My Spanish teacher asked me to turn in my essay,30
post,3jrus0,2qh72,jokes,false,1441479449,https://old.reddit.com/r/Jokes/comments/3jrus0/dog_for_sale/,self.jokes,,Eats everything. Loves kids.,Dog for sale,2
post,3jruor,2qh72,jokes,false,1441479404,https://old.reddit.com/r/Jokes/comments/3jruor/whats_the_difference_between_a_beta_a_worm_and_a/,self.jokes,,[deleted],"what's the difference between a beta, a worm, and a patient with dementia?",0
post,3jrulo,2qh72,jokes,false,1441479367,https://old.reddit.com/r/Jokes/comments/3jrulo/sir_there_is_a_complaint_filed_against_you_you/,self.jokes,,"OK. Who filed the complaint, prime minister or the whore?","Sir, there is a complaint filed against you. You called the prime minister a whore...",0
post,3jrsrz,2qh72,jokes,false,1441478529,https://old.reddit.com/r/Jokes/comments/3jrsrz/garry_glitter_gave_me_my_first_guitar_lesson_the/,self.jokes,,He showed me how to finger A minor ,Garry Glitter gave me my first guitar lesson the other day,7
post,3jrsnz,2qh72,jokes,false,1441478479,https://old.reddit.com/r/Jokes/comments/3jrsnz/make_a_sentence_with_the_following_words_elephant/,self.jokes,,Ant in an elephant's ass,Make a sentence with the following words 'elephant' 'ant' 'ass' 'in' and 'bamboo',0
post,3jrsjm,2qh72,jokes,false,1441478427,https://old.reddit.com/r/Jokes/comments/3jrsjm/did_you_hear_about_the_clairvoyant_midget_that/,self.jokes,,He's a small medium at large.,Did you hear about the clairvoyant midget that escaped from jail?,11
post,3jrsfe,2qh72,jokes,false,1441478368,https://old.reddit.com/r/Jokes/comments/3jrsfe/i_started_crossfit_yesterday/,self.jokes,,And my throat is killing me,I started crossfit yesterday,2
post,3jrrf5,2qh72,jokes,false,1441477882,https://old.reddit.com/r/Jokes/comments/3jrrf5/a_dyslexic_agnostic_insomniac/,self.jokes,,"A dyslexic, agnostic insomniac lay awake all night wondering if there is a dog. 

EDIT: Credit to David Foster Wallace. ","A dyslexic, agnostic insomniac",38
post,3jrrbp,2qh72,jokes,false,1441477842,https://old.reddit.com/r/Jokes/comments/3jrrbp/midget_with_a_speech_impediment/,self.jokes,,"A guy calls a horse rancher and says he’s sending a friend over to look at a race horse he wants to buy. 
The rancher says “how will I recognize him?” 
""Easy, he’s a midget with a speech impediment”
The midget shows up and the rancher asks him if he is looking for a male or female horse. 
""A female horth” So he shows him a prized filly. 
""Nith lookin’ horth. Can I thee her eyeth?"" 
So the rancher picks up the midget and gets him eye to eye with the horse. Puts him down. 
""Nith eyeth, can I thee her earzth?” 
The rancher picks up the little fella again and shows him the horse’s ears. Puts him down. 
""Hmm, nith earzth. Can I thee her mouf?” The rancher is getting impatient with having to lift the midget every time he asks a question, but he picks him up again and shows him the horse’s mouth. ""Hmm, nith mouf, can I thee her twat?” Totally pissed off at this point, the rancher grabs him under his arm and jams the midget’s head as far as he can up the horse’s twat, pulls him out and slams him on the ground.
The midget gets up, sputtering and coughing and says, “Perhapth, I should rephrathe that. Can I thee her wun awound a widdle bit?”",Midget with a speech impediment.,82
post,3jrr9u,2qh72,jokes,false,1441477816,https://old.reddit.com/r/Jokes/comments/3jrr9u/you_know_what_the_number_one_leading_cause_of/,self.jokes,,"Sexy kids.

(Pro Tip: I tell this to every single one of my First Dates. It's my Late 20s testing threshold for whether or not they'll tolerate me for very long.)

Edit: and no, I don't mean them tolerating my proclivity toward sexy kids.

Edit2: and no, I don't see any kids as being sexy.

Edit3: except some of the Disney Channel stars from a decade-plus-ago, when I was a teenager, too. And it's kind of trippy to see those old episodes now and you're time traveling inside your head, like you're that age again. And you're able to remember what made them attractive to you. That's a mind-fuck.

Edit4: How did my last date go? It went alright. We fucked all night then I told her the joke since I was afraid it would scare her away like the last few girls, and I was feeling lonely lately. We were both tired, naked, and sweaty. I told her the joke. She laughed but said, ""That's atrocious!"" And I said, ""That's a mighty big word for a twelve year old.""

Edit5: I'll be here all week.

Edit6: I'll be incarcerated next week.

Edit7: confession time: I ripped this joke off my pastor. It was payback for him ripping off my clothes.

Edit8: that last edit wasn't a joke. My pastor ruined perfectly good clothes my mom purchased for me every Christmas. Sunday masses were a bummer cause I got all dressed up and he couldn't control himself. It's tough being young and wanting to be fashionable. It's my fault. My ass looked good in those jeans.

Edit9: for anyone who thinks I'm making light of pedophilia, it's okay. I'm allowed to. I have plenty of pedophile friends.

Edit10: my boss at my first job was right about networking. My name isn't Jared for nothing.

Edit11: but seriously, go visit victimsofcrime DOT org if you know of anyone currently in a crisis. You could be seriously saving someone from a life of therapy and self-torture. Thank you for laughing, if you did. And thank you for reading this far, at least, if you didn't laugh. I gotta go now. This cop has been staring me down all morning. Can't a single guy watch kids play at the park in peace? Geez.

Edit12: apparently, some of you think this joke has too many edits. I guess I should have posted to to /r/TrueJokes instead.

Edit13: spellcheck 

Edit14: omgfrontpage and guilded. Wow, first post, too. Wow. Thank you. I'm gonna go touch a child a child for every upvote I get.

Edit15: this whole post is becoming stale. It's like beating off on a dead child.","You know what the number one leading cause of pedophilia is, right?",17
post,3jrqya,2qh72,jokes,false,1441477679,https://old.reddit.com/r/Jokes/comments/3jrqya/did_you_hear_about_the_two_jamaican_turtles_at/,self.jokes,,They were just looking for Michelle Bachman. ,Did you hear about the two Jamaican Turtles at the RNC?,2
post,3jrpyv,2qh72,jokes,false,1441477262,https://old.reddit.com/r/Jokes/comments/3jrpyv/dad_jokes_for_fathers_day/,self.jokes,,"Hey guys! It's father's day in Australia today, so how about your best, most eye-rollingest guffaw-inducing dad jokes? Hit me with your best shot!",Dad jokes for Father's day,0
post,3jrpea,2qh72,jokes,false,1441476996,https://old.reddit.com/r/Jokes/comments/3jrpea/what_do_you_call_a_football_team_full_of_retards/,self.jokes,,Special teams.,What do you call a football team full of retards?,2
post,3jrpa4,2qh72,jokes,false,1441476944,https://old.reddit.com/r/Jokes/comments/3jrpa4/american_politics/,self.jokes,,[deleted],American Politics,6
post,3jrp2z,2qh72,jokes,false,1441476857,https://old.reddit.com/r/Jokes/comments/3jrp2z/what_comes_between_fear_and_sex/,self.jokes,,Fünf,What comes between fear and sex?,11
post,3jrnyf,2qh72,jokes,false,1441476315,https://old.reddit.com/r/Jokes/comments/3jrnyf/a_group_of_guys_all_aged_about_40_discussed_where/,self.jokes,,"Finally it was agreed that they would meet at the Ocean View restaurant because the waitresses there were pretty.

Ten years later, at age 50, the friends once again discussed where they should meet for lunch.Finally it was agreed that they would meet at the Ocean View restaurant because the food was good and the wine selection was excellent.


Ten years later, at age 60, the friends again discussed where they should meet for lunch.Finally it was agreed that they would meet at the Ocean View restaurant because they could dine in peace and quiet and the restaurant had a beautiful view of the ocean.

Ten years later, at age 70, the friends discussed where they should meet for lunch.
Finally it was agreed that they would meet at the Ocean View restaurant because the restaurant was wheelchair accessible and had an elevator.

Ten years later, at age 80, the friends discussed where they should meet for lunch.
Finally it was agreed that they would meet at the Ocean View restaurant because they had never been there before.","A group of guys, all aged about 40, discussed where they should meet for lunch",720
post,3jrnlp,2qh72,jokes,false,1441476150,https://old.reddit.com/r/Jokes/comments/3jrnlp/dont_eat_the_vegetables_in_hospital_cafeterias/,self.jokes,,"The police track you down after that, you see.",Don't eat the vegetables in hospital cafeterias,3
post,3jrmoc,2qh72,jokes,false,1441475730,https://old.reddit.com/r/Jokes/comments/3jrmoc/whats_the_best_part_about_fucking_21_year_olds/,self.jokes,,[deleted],What's the best part about fucking 21 year olds?,0
post,3jrmfj,2qh72,jokes,false,1441475609,https://old.reddit.com/r/Jokes/comments/3jrmfj/whats_a_cats_favorite_song/,self.jokes,,3 blind mice,What's a cats favorite song?,0
post,3jrmb2,2qh72,jokes,false,1441475552,https://old.reddit.com/r/Jokes/comments/3jrmb2/are_youre_hungry_now/,self.jokes,,Cause I'm Hungarian!,Are you're hungry now?,0
post,3jrm13,2qh72,jokes,false,1441475430,https://old.reddit.com/r/Jokes/comments/3jrm13/what_do_you_call_a_man_whos_on_fire/,self.jokes,,Bernie. ,What do you call a man who's on fire?,0
post,3jrljn,2qh72,jokes,false,1441475181,https://old.reddit.com/r/Jokes/comments/3jrljn/an_angel_and_a_man/,self.jokes,,"An angel appears in a puff of smoke to a man and says to him, ""Because you have lived a good and virtuous life, I can offer you a gift: you can be the most handsome man in the world, or you can have infinite wisdom, or you can have limitless wealth.""
Reflecting on his life, the man says, ""I'll take the wisdom.""
""Wisdom is yours,"" says the angel, disappearing in another puff.
The smoke is barely clear before the man thinks, ""I should have taken the money.""",An angel and a man,320
post,3jrkvx,2qh72,jokes,false,1441474877,https://old.reddit.com/r/Jokes/comments/3jrkvx/try_saying_i_heaven_this_order_three_times/,self.jokes,,Nothing wrong if you do :),"Try saying ""I heaven this order"" three times.",0
post,3jrkvk,2qh72,jokes,false,1441474873,https://old.reddit.com/r/Jokes/comments/3jrkvk/what_did_the_third_reich_say_when_they_fired/,self.jokes,,"""You're ladolf.""",What did the Third Reich say when they fired Hitler?,0
post,3jrkkc,2qh72,jokes,false,1441474724,https://old.reddit.com/r/Jokes/comments/3jrkkc/if_youd_like_to_know_whats_in_style_right_now/,self.jokes,,I've heard shirts with collars are really poppin.,If you'd like to know what's in style right now...,0
post,3jrj7q,2qh72,jokes,false,1441474099,https://old.reddit.com/r/Jokes/comments/3jrj7q/two_blonde_girls_are_heading_to_disneyland/,self.jokes,,"While driving they see a sign ""Disney Left"". They cry and head home.

(Little bro told me this one. Not sure if it has been told before.)",Two blonde girls are heading to Disneyland...,6
post,3jrin9,2qh72,jokes,false,1441473828,https://old.reddit.com/r/Jokes/comments/3jrin9/how_does_the_mummy_plan_to_destroy_superman/,self.jokes,,He's going to lure him into the crypt tonight.,How does the mummy plan to destroy Superman?,90
post,3jril4,2qh72,jokes,false,1441473802,https://old.reddit.com/r/Jokes/comments/3jril4/sex_vs_frisbee/,self.jokes,,"Casual sex is like playing Frisbee. It's not something I think about doing all the time but if the opportunity presents itself and you have the time it's hard to justify saying no. It's usually fun. Sometimes it sucks because your timing is off,you try some fancy moves that made perfect sense in your head but not so much in execution,the other person can't throw or you get something in your eye. But for the most part its fun. Everyone walks away smiling and when you remember it you think, that was a good time. I should do that more often.
If you read this and think I'm totally off base consider this: 1.you don't like frisbee 2.you have never played frisbee with someone that was good at it. 3.your perception of frisbee is not really frisbee. It's golf.",Sex vs Frisbee,3
post,3jri1y,2qh72,jokes,false,1441473547,https://old.reddit.com/r/Jokes/comments/3jri1y/erections_happen_all_the_time/,self.jokes,,"A man is about to get a prostate exam from his doctor. Before the doctor begins, he tells the man ""I must tell you, during this type of examination, erections happen all the time. They are very common, and trust me, it's nothing to be embarrassed about.""

The man seems a little uncomfortable, but the doctor continues, ""Now a little less common, is you may get one too.""",Erections happen all the time,444
post,3jrh6k,2qh72,jokes,false,1441473145,https://old.reddit.com/r/Jokes/comments/3jrh6k/two_murcians_in_a_bar_talk_about_the_refugee/,self.jokes,,"Dude what's your thought about those refugees?

I dunno, but Europeans need to something before it's too late!

Native American joins in: Yep, we completely underestimated them.",Two Murcians in a bar talk about the refugee crisis,2
post,3jrh69,2qh72,jokes,false,1441473141,https://old.reddit.com/r/Jokes/comments/3jrh69/how_do_you_spot_an_attention_whore_on_reddit/,self.jokes,,[-],How do you spot an attention whore on reddit?,0
post,3jrh2c,2qh72,jokes,false,1441473095,https://old.reddit.com/r/Jokes/comments/3jrh2c/what_do_you_call/,self.jokes,,"What do you call nuts on a wall?
Walnuts
What do you call nuts on a chest? 
Chestnuts
What do you call nuts on a chin?
A dick in the mouth ",What do you call?,2
post,3jrgbj,2qh72,jokes,false,1441472751,https://old.reddit.com/r/Jokes/comments/3jrgbj/i_met_mike_tyson_and_he_had_his_tiger_with_him_i/,self.jokes,,"He said, ""Well you were mythtaken.""","I met Mike Tyson and he had his tiger with him. I said, ""Wow! I can't believe you actually have a tiger! I thought that was a myth.""",67
post,3jrf4n,2qh72,jokes,false,1441472196,https://old.reddit.com/r/Jokes/comments/3jrf4n/how_come_dinosaurs_dont_talk/,self.jokes,,[deleted],How come dinosaurs don't talk?,0
post,3jren6,2qh72,jokes,false,1441471958,https://old.reddit.com/r/Jokes/comments/3jren6/what_is_six_inches_long_has_a_bald_head_and/,self.jokes,,100$ bill,What is six inches long has a bald head and drives every woman crazy?,1
post,3jrehq,2qh72,jokes,false,1441471893,https://old.reddit.com/r/Jokes/comments/3jrehq/whats_red_bloody_and_hangs_of_the_back_of_a_train/,self.jokes,,Miscarriage.,"What's red, bloody and hangs of the back of a train?",0
post,3jree3,2qh72,jokes,false,1441471846,https://old.reddit.com/r/Jokes/comments/3jree3/two_jihadis_walked_in_to_a_bar/,self.jokes,,They didn't blow it up. ,Two Jihadis Walked In to a bar,1
post,3jrdpj,2qh72,jokes,false,1441471525,https://old.reddit.com/r/Jokes/comments/3jrdpj/what_did_the_premature_ejaculatist_say_to_his/,self.jokes,,"Sorry... 


That came out wrong.",What did the premature ejaculatist say to his offended lover?,21
post,3jrdp0,2qh72,jokes,false,1441471516,https://old.reddit.com/r/Jokes/comments/3jrdp0/a_man_goes_to_the_doctor_he_says_hes_depressed/,self.jokes,,"The man bursts into tears and replies: but, Doctor... I *am* Pagliacci.","A man goes to the Doctor. He says he's depressed. Life seems harsh, cruel, and what lies ahead is vague and uncertain. The Doctor says: The treatment's simple, a great clown named Pagliacci is in town, go and see him! That should pick you up.",1
post,3jrda4,2qh72,jokes,false,1441471335,https://old.reddit.com/r/Jokes/comments/3jrda4/taking_the_lives_away_from_12_baby_chicks/,self.jokes,,Bought an egg carton at the grocery store...,Taking the lives away from 12 baby chicks.,0
post,3jrcuw,2qh72,jokes,false,1441471125,https://old.reddit.com/r/Jokes/comments/3jrcuw/two_couples_were_playing_cards_john_accidentally/,self.jokes,,"Two couples were playing cards. John accidentally dropped some cards on the floor. When he bent down under the table to pick them up, he noticed .... Bill's wife was not wearing any panties! Shocked by this, John hit his head on the table and emerged red-faced.

Later, John went to the kitchen to get some refreshments. Bill's wife followed him and asked, ""Did you see anything that you liked under there?""

John admitted that, well, yes he did.

She said ""You can have it, but it will cost you $100.""

After a minute or two, John indicates that he is interested. She tells him that since Bill works Friday afternoons and John doesn't, John should come to her house around 2:00 p.m. on Friday.

Friday came and John went to her house at 2:00 p.m. After paying her $100 they went to the bedroom, had sex, and then John left.

Bill came home about 6:00 P.M. He asked his wife, ""Did John come by this afternoon?""

Reluctantly, she replied, ""Yes, he did stop by for a few minutes.""

Next Bill asked, ""Did John give you $100?""

She thinks 'Oh hell, he knows!' Finally she says, ""Yes, he did give me $100.""

""Good,"" Bill says. ""John came by the office this morning and borrowed $100 from me. He said that he would stop by our house on his way home and pay me back.","Two couples were playing cards. John accidentally dropped some cards on the floor. When he bent down under the table to pick them up, he noticed....",3934
post,3jrcmt,2qh72,jokes,false,1441471025,https://old.reddit.com/r/Jokes/comments/3jrcmt/when_will_the_jared_jokes_stop/,self.jokes,,When they get too old.,When will the Jared jokes stop?,215
post,3jrcmb,2qh72,jokes,false,1441471022,https://old.reddit.com/r/Jokes/comments/3jrcmb/facebook_keeps_me_from_talking_to_people/,self.jokes,,[deleted],Facebook keeps me from talking to people,0
post,3jrbuv,2qh72,jokes,false,1441470660,https://old.reddit.com/r/Jokes/comments/3jrbuv/we_all_know_what_this_means/,self.jokes,,"🎺🎺🎺🎺



It's just 4 trumpets! 
Or ITS JOHN CENA 

🎺🎺🎺🎺
Sorry.",We all know what this means,0
post,3jrbr1,2qh72,jokes,false,1441470607,https://old.reddit.com/r/Jokes/comments/3jrbr1/i_am_here_folks/,self.jokes,,[removed],I am here folks,0
post,3jr7iu,2qh72,jokes,false,1441468668,https://old.reddit.com/r/Jokes/comments/3jr7iu/noahs_diary_day_39/,self.jokes,,[deleted],Noah's diary day 39,73
post,3jr7eo,2qh72,jokes,false,1441468611,https://old.reddit.com/r/Jokes/comments/3jr7eo/a_dyslexic_walks_into_a_bra/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jr7eo/a_dyslexic_walks_into_a_bra/,,A dyslexic walks into a bra...,1
post,3jr74v,2qh72,jokes,false,1441468483,https://old.reddit.com/r/Jokes/comments/3jr74v/knock_knock/,self.jokes,,[deleted],"Knock, Knock...",1
post,3jr60g,2qh72,jokes,false,1441467965,https://old.reddit.com/r/Jokes/comments/3jr60g/how_do_you_spot_an_attention_whore_on_reddit/,self.jokes,,"Edit: Wow, I did not expect this to get so many upvotes!",How do you spot an attention whore on reddit?,0
post,3jr5sq,2qh72,jokes,false,1441467871,https://old.reddit.com/r/Jokes/comments/3jr5sq/a_man_with_a_stutter/,self.jokes,,"A man with a stutter is visiting the doctor.

""How's the stutter?"", asks the doctor.

""It's g-getting better. My mate calls me D-Donkey,"" replies the man.

""Any idea why?"" The doctor asks.

""No, but he aw he aw he aw he always calls me that.""",A man with a stutter...,620
post,3jr585,2qh72,jokes,false,1441467623,https://old.reddit.com/r/Jokes/comments/3jr585/whats_the_difference_between_a_viola_and_a_bouncy/,self.jokes,,"You take your shoes off to jump on a bouncy castle.

(From a guitarist/pianist/bass/banjo/mandolin player friend who despises classical instruments.)",What's the difference between a Viola and a Bouncy Castle.,0
post,3jr4dc,2qh72,jokes,false,1441467253,https://old.reddit.com/r/Jokes/comments/3jr4dc/why_does_michael_j_fox_make_the_best_milkshakes/,self.jokes,,Because he only uses the finest ingredients. ,Why does Michael J Fox make the best milkshakes?,4
post,3jr43h,2qh72,jokes,false,1441467135,https://old.reddit.com/r/Jokes/comments/3jr43h/help/,self.jokes,,I can't post anything on Reddit! Pls help!,Help!,0
post,3jr41x,2qh72,jokes,false,1441467114,https://old.reddit.com/r/Jokes/comments/3jr41x/if_i_told_you_you_have_a_beautiful_body/,self.jokes,,would you hold it against me?,if i told you you have a beautiful body....,0
post,3jr406,2qh72,jokes,false,1441467090,https://old.reddit.com/r/Jokes/comments/3jr406/françois_hollande/,self.jokes,https://www.reddit.com/r/Jokes/comments/3jr406/françois_hollande/,,François Hollande.,3
post,3jr3ms,2qh72,jokes,false,1441466920,https://old.reddit.com/r/Jokes/comments/3jr3ms/a_crusty_old_sergeant_major_walks_into_a_brothel/,self.jokes,,"He walks up to the receptionist and says, ""I'm a sergeant major, I've seen combat in every major conflict for the last 35 years, and I want the best goddamn hooker you've got in this place!""

The receptionist nods and leads him to one of the back rooms. Waiting there is a stunningly beautiful woman. The sergeant major  tells the receptionist to leave and starts making small talk with the hooker.

""So,"" the hooker says. ""What makes you worth my time?""

The sergeant major replies, ""I'm a goddamn sergeant major and I've seen combat in every conflict in the last 35 years! I wear command presence like you wear a skimpy skirt, and I'll prove it to you!"" The sergeant major takes off his pants, looks down at his penis, and says, ""Dick! Atten-SHUN!"" His manlihood instantly snaps to the position of attention.

The hooker's eyes get wide. ""That's incredible!""

""Yes,"" the sergeant major says. ""It is. Now, watch this."" He looks back down, and says ""At ease!"" His member returns to its flaccid state.

The hooker is, again, impressed. She asks if he can do it again, and he does. Twice. Finally, she says, ""Well, let's get to it, shall we?""

The sergeant major, just for good measure, looks down and says, ""Dick! Atten-SHUN!"" one more time. But this time, nothing happens. The sergeant major growls in anger.

""Dick! Atten-SHUN!"" Still, nothing happens.

The sergeant major jumps over into the corner and starts vigorously beating his meat.

""What are you doing?!"" the hooker exclaims.

""This little soldier won't listen to me!"" the sergeant major shouts, ""So I'm giving him a dishonorable discharge!""",A crusty old sergeant major walks into a brothel in Korea...,111
post,3jr3mb,2qh72,jokes,false,1441466914,https://old.reddit.com/r/Jokes/comments/3jr3mb/what_the_difference_between_a_violin_and_a_viola/,self.jokes,,[deleted],What the difference between a Violin and a Viola?,0
post,3jr3dd,2qh72,jokes,false,1441466802,https://old.reddit.com/r/Jokes/comments/3jr3dd/i_tried_taking_a_shower_while_my_water_softener/,self.jokes,,[deleted],"I tried taking a shower while my water softener was broken, but it was hard",1
post,3jr3br,2qh72,jokes,false,1441466782,https://old.reddit.com/r/Jokes/comments/3jr3br/why_didnt_isaac_newton_drink_wine/,self.jokes,,He knew better than to drink and derive.,Why didn't Isaac Newton drink wine?,38
post,3jr2t9,2qh72,jokes,false,1441466521,https://old.reddit.com/r/Jokes/comments/3jr2t9/life_as_a_drunk_has_never_been_easy/,self.jokes,,[deleted],Life as a drunk has never been easy,0
post,3jr2t7,2qh72,jokes,false,1441466521,https://old.reddit.com/r/Jokes/comments/3jr2t7/why_isnt_sean_connery_allowed_to_play_super_mario/,self.jokes,,He kept trying to shave the princess.,Why isn't Sean Connery allowed to play Super Mario Bros. any more?,18
post,3jr1zz,2qh72,jokes,false,1441466116,https://old.reddit.com/r/Jokes/comments/3jr1zz/went_to_the_store_to_buy_some_condoms/,self.jokes,,[deleted],Went to the Store to buy some Condoms,0
post,3jr1l4,2qh72,jokes,false,1441465904,https://old.reddit.com/r/Jokes/comments/3jr1l4/kids_say_the_darnedest_things/,self.jokes,,"A young lad was in the car with his Dad on the way home. Dad's listening to the radio to hear the football scores. They get stopped by a routine police patrol who do a quick licence check and send them on their way. Flummoxed by this, the boy asks his father who those people were. Not listening, the father says, ""bastards"" (as he's just heard his favourite team have lost 1-0). Arriving home they wipe their feet on the welcome mat. Dad drops his keys and exclaims, ""Shite!"". The boy walks into the house and heads to the kitchen while his father goes upstairs. ""Mammy, what are you doing?"", he asks as he a